-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jan 11 2025 14:15:47

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MMU" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MMU
entity MMU is
port (
    ORA : out std_logic_vector(7 downto 0);
    A : in std_logic_vector(15 downto 0);
    CXXXOUT : out std_logic;
    ROMEN1_N : inout std_logic;
    Q3 : in std_logic;
    R_W_N_245 : inout std_logic;
    ROMEN2_N : out std_logic;
    INH_N : in std_logic;
    EN80_N : out std_logic;
    DMA_N : in std_logic;
    MD7 : inout std_logic;
    CASEN_N : out std_logic;
    KBD_N : out std_logic;
    R_W_N : in std_logic;
    PRAS_N : in std_logic;
    PHI_0 : in std_logic);
end MMU;

-- Architecture of MMU
-- View name is \INTERFACE\
architecture \INTERFACE\ of MMU is

signal \N__6167\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6138\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5595\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5382\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5376\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5364\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5046\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4605\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4503\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4222\ : std_logic;
signal \N__4219\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4158\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4030\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4012\ : std_logic;
signal \N__4009\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3991\ : std_logic;
signal \N__3988\ : std_logic;
signal \N__3985\ : std_logic;
signal \N__3984\ : std_logic;
signal \N__3981\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3975\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3949\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3933\ : std_logic;
signal \N__3930\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3921\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3907\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3870\ : std_logic;
signal \N__3867\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3858\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3852\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3821\ : std_logic;
signal \N__3818\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3809\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3799\ : std_logic;
signal \N__3796\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3787\ : std_logic;
signal \N__3784\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3751\ : std_logic;
signal \N__3748\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3714\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3693\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3687\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3679\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3655\ : std_logic;
signal \N__3654\ : std_logic;
signal \N__3651\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3603\ : std_logic;
signal \N__3602\ : std_logic;
signal \N__3599\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3593\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3582\ : std_logic;
signal \N__3579\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3575\ : std_logic;
signal \N__3570\ : std_logic;
signal \N__3567\ : std_logic;
signal \N__3564\ : std_logic;
signal \N__3561\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3550\ : std_logic;
signal \N__3545\ : std_logic;
signal \N__3542\ : std_logic;
signal \N__3539\ : std_logic;
signal \N__3536\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3530\ : std_logic;
signal \N__3527\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3525\ : std_logic;
signal \N__3524\ : std_logic;
signal \N__3521\ : std_logic;
signal \N__3518\ : std_logic;
signal \N__3517\ : std_logic;
signal \N__3514\ : std_logic;
signal \N__3511\ : std_logic;
signal \N__3510\ : std_logic;
signal \N__3505\ : std_logic;
signal \N__3502\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3491\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3479\ : std_logic;
signal \N__3476\ : std_logic;
signal \N__3473\ : std_logic;
signal \N__3470\ : std_logic;
signal \N__3467\ : std_logic;
signal \N__3464\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3460\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3452\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3446\ : std_logic;
signal \N__3443\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3437\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3428\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3419\ : std_logic;
signal \N__3416\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3411\ : std_logic;
signal \N__3410\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3403\ : std_logic;
signal \N__3398\ : std_logic;
signal \N__3395\ : std_logic;
signal \N__3392\ : std_logic;
signal \N__3391\ : std_logic;
signal \N__3388\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3382\ : std_logic;
signal \N__3379\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3377\ : std_logic;
signal \N__3376\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3372\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3361\ : std_logic;
signal \N__3354\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3345\ : std_logic;
signal \N__3342\ : std_logic;
signal \N__3335\ : std_logic;
signal \N__3332\ : std_logic;
signal \N__3323\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3314\ : std_logic;
signal \N__3311\ : std_logic;
signal \N__3308\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3298\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3295\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3293\ : std_logic;
signal \N__3292\ : std_logic;
signal \N__3275\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3266\ : std_logic;
signal \N__3263\ : std_logic;
signal \N__3260\ : std_logic;
signal \N__3257\ : std_logic;
signal \N__3254\ : std_logic;
signal \N__3251\ : std_logic;
signal \N__3248\ : std_logic;
signal \N__3245\ : std_logic;
signal \N__3242\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3236\ : std_logic;
signal \N__3235\ : std_logic;
signal \N__3232\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3229\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3208\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3200\ : std_logic;
signal \N__3197\ : std_logic;
signal \N__3194\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3177\ : std_logic;
signal \N__3170\ : std_logic;
signal \N__3167\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3163\ : std_logic;
signal \N__3162\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3157\ : std_logic;
signal \N__3152\ : std_logic;
signal \N__3147\ : std_logic;
signal \N__3146\ : std_logic;
signal \N__3141\ : std_logic;
signal \N__3138\ : std_logic;
signal \N__3135\ : std_logic;
signal \N__3132\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3122\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3103\ : std_logic;
signal \N__3100\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3094\ : std_logic;
signal \N__3089\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3083\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3077\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3071\ : std_logic;
signal \N__3068\ : std_logic;
signal \N__3065\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3058\ : std_logic;
signal \N__3055\ : std_logic;
signal \N__3052\ : std_logic;
signal \N__3051\ : std_logic;
signal \N__3048\ : std_logic;
signal \N__3045\ : std_logic;
signal \N__3042\ : std_logic;
signal \N__3035\ : std_logic;
signal \N__3032\ : std_logic;
signal \N__3029\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3022\ : std_logic;
signal \N__3019\ : std_logic;
signal \N__3016\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3005\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2996\ : std_logic;
signal \N__2993\ : std_logic;
signal \N__2990\ : std_logic;
signal \N__2987\ : std_logic;
signal \N__2984\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2978\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2962\ : std_logic;
signal \N__2961\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2950\ : std_logic;
signal \N__2949\ : std_logic;
signal \N__2948\ : std_logic;
signal \N__2945\ : std_logic;
signal \N__2942\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2927\ : std_logic;
signal \N__2924\ : std_logic;
signal \N__2921\ : std_logic;
signal \N__2918\ : std_logic;
signal \N__2915\ : std_logic;
signal \N__2912\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2906\ : std_logic;
signal \N__2903\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2890\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2882\ : std_logic;
signal \N__2879\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2873\ : std_logic;
signal \N__2870\ : std_logic;
signal \N__2867\ : std_logic;
signal \N__2864\ : std_logic;
signal \N__2861\ : std_logic;
signal \N__2858\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2846\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2837\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2833\ : std_logic;
signal \N__2830\ : std_logic;
signal \N__2827\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2816\ : std_logic;
signal \N__2813\ : std_logic;
signal \N__2812\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2808\ : std_logic;
signal \N__2805\ : std_logic;
signal \N__2802\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2794\ : std_logic;
signal \N__2791\ : std_logic;
signal \N__2788\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2780\ : std_logic;
signal \N__2777\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2768\ : std_logic;
signal \N__2765\ : std_logic;
signal \N__2762\ : std_logic;
signal \N__2759\ : std_logic;
signal \N__2756\ : std_logic;
signal \N__2753\ : std_logic;
signal \N__2750\ : std_logic;
signal \N__2747\ : std_logic;
signal \N__2744\ : std_logic;
signal \N__2741\ : std_logic;
signal \N__2738\ : std_logic;
signal \N__2735\ : std_logic;
signal \N__2732\ : std_logic;
signal \N__2729\ : std_logic;
signal \N__2726\ : std_logic;
signal \N__2723\ : std_logic;
signal \N__2720\ : std_logic;
signal \N__2717\ : std_logic;
signal \N__2714\ : std_logic;
signal \N__2711\ : std_logic;
signal \N__2708\ : std_logic;
signal \N__2707\ : std_logic;
signal \N__2702\ : std_logic;
signal \N__2701\ : std_logic;
signal \N__2698\ : std_logic;
signal \N__2695\ : std_logic;
signal \N__2690\ : std_logic;
signal \N__2687\ : std_logic;
signal \N__2684\ : std_logic;
signal \N__2681\ : std_logic;
signal \N__2678\ : std_logic;
signal \N__2675\ : std_logic;
signal \N__2672\ : std_logic;
signal \N__2671\ : std_logic;
signal \N__2670\ : std_logic;
signal \N__2665\ : std_logic;
signal \N__2662\ : std_logic;
signal \N__2657\ : std_logic;
signal \N__2654\ : std_logic;
signal \N__2651\ : std_logic;
signal \N__2648\ : std_logic;
signal \N__2645\ : std_logic;
signal \N__2642\ : std_logic;
signal \N__2639\ : std_logic;
signal \N__2636\ : std_logic;
signal \N__2633\ : std_logic;
signal \N__2630\ : std_logic;
signal \N__2627\ : std_logic;
signal \N__2624\ : std_logic;
signal \N__2621\ : std_logic;
signal \N__2618\ : std_logic;
signal \N__2615\ : std_logic;
signal \N__2612\ : std_logic;
signal \N__2609\ : std_logic;
signal \N__2606\ : std_logic;
signal \N__2603\ : std_logic;
signal \N__2600\ : std_logic;
signal \N__2597\ : std_logic;
signal \N__2594\ : std_logic;
signal \N__2591\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2585\ : std_logic;
signal \N__2584\ : std_logic;
signal \N__2581\ : std_logic;
signal \N__2578\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2572\ : std_logic;
signal \N__2569\ : std_logic;
signal \N__2564\ : std_logic;
signal \N__2561\ : std_logic;
signal \N__2558\ : std_logic;
signal \N__2555\ : std_logic;
signal \N__2552\ : std_logic;
signal \N__2549\ : std_logic;
signal \N__2548\ : std_logic;
signal \N__2545\ : std_logic;
signal \N__2542\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2536\ : std_logic;
signal \N__2533\ : std_logic;
signal \N__2530\ : std_logic;
signal \N__2525\ : std_logic;
signal \N__2522\ : std_logic;
signal \N__2519\ : std_logic;
signal \N__2518\ : std_logic;
signal \N__2515\ : std_logic;
signal \N__2512\ : std_logic;
signal \N__2511\ : std_logic;
signal \N__2508\ : std_logic;
signal \N__2505\ : std_logic;
signal \N__2502\ : std_logic;
signal \N__2499\ : std_logic;
signal \N__2492\ : std_logic;
signal \N__2489\ : std_logic;
signal \N__2486\ : std_logic;
signal \N__2483\ : std_logic;
signal \N__2480\ : std_logic;
signal \N__2477\ : std_logic;
signal \N__2474\ : std_logic;
signal \N__2471\ : std_logic;
signal \N__2468\ : std_logic;
signal \N__2465\ : std_logic;
signal \N__2462\ : std_logic;
signal \N__2459\ : std_logic;
signal \N__2456\ : std_logic;
signal \N__2453\ : std_logic;
signal \N__2450\ : std_logic;
signal \N__2447\ : std_logic;
signal \N__2444\ : std_logic;
signal \N__2441\ : std_logic;
signal \N__2438\ : std_logic;
signal \N__2437\ : std_logic;
signal \N__2436\ : std_logic;
signal \N__2435\ : std_logic;
signal \N__2430\ : std_logic;
signal \N__2427\ : std_logic;
signal \N__2424\ : std_logic;
signal \N__2421\ : std_logic;
signal \N__2418\ : std_logic;
signal \N__2415\ : std_logic;
signal \N__2412\ : std_logic;
signal \N__2407\ : std_logic;
signal \N__2404\ : std_logic;
signal \N__2401\ : std_logic;
signal \N__2396\ : std_logic;
signal \N__2393\ : std_logic;
signal \N__2390\ : std_logic;
signal \N__2389\ : std_logic;
signal \N__2386\ : std_logic;
signal \N__2383\ : std_logic;
signal \N__2378\ : std_logic;
signal \N__2375\ : std_logic;
signal \N__2372\ : std_logic;
signal \N__2369\ : std_logic;
signal \N__2366\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2360\ : std_logic;
signal \N__2357\ : std_logic;
signal \N__2356\ : std_logic;
signal \N__2353\ : std_logic;
signal \N__2350\ : std_logic;
signal \N__2345\ : std_logic;
signal \N__2342\ : std_logic;
signal \N__2339\ : std_logic;
signal \N__2336\ : std_logic;
signal \N__2333\ : std_logic;
signal \N__2330\ : std_logic;
signal \N__2327\ : std_logic;
signal \N__2324\ : std_logic;
signal \N__2321\ : std_logic;
signal \N__2318\ : std_logic;
signal \N__2317\ : std_logic;
signal \N__2314\ : std_logic;
signal \N__2311\ : std_logic;
signal \N__2306\ : std_logic;
signal \N__2303\ : std_logic;
signal \N__2300\ : std_logic;
signal \N__2299\ : std_logic;
signal \N__2298\ : std_logic;
signal \N__2295\ : std_logic;
signal \N__2292\ : std_logic;
signal \N__2289\ : std_logic;
signal \N__2282\ : std_logic;
signal \N__2279\ : std_logic;
signal \N__2276\ : std_logic;
signal \N__2273\ : std_logic;
signal \N__2270\ : std_logic;
signal \N__2267\ : std_logic;
signal \N__2264\ : std_logic;
signal \N__2261\ : std_logic;
signal \N__2258\ : std_logic;
signal \N__2255\ : std_logic;
signal \N__2252\ : std_logic;
signal \N__2249\ : std_logic;
signal \N__2246\ : std_logic;
signal \N__2243\ : std_logic;
signal \N__2240\ : std_logic;
signal \N__2237\ : std_logic;
signal \N__2234\ : std_logic;
signal \N__2231\ : std_logic;
signal \N__2228\ : std_logic;
signal \N__2225\ : std_logic;
signal \N__2222\ : std_logic;
signal \N__2219\ : std_logic;
signal \N__2216\ : std_logic;
signal \N__2213\ : std_logic;
signal \N__2210\ : std_logic;
signal \N__2207\ : std_logic;
signal \N__2204\ : std_logic;
signal \N__2201\ : std_logic;
signal \N__2198\ : std_logic;
signal \N__2197\ : std_logic;
signal \N__2194\ : std_logic;
signal \N__2191\ : std_logic;
signal \N__2186\ : std_logic;
signal \N__2183\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U_R_W_N_245LegalizeSB_DFFNet\ : std_logic;
signal \DMA_N_c\ : std_logic;
signal \R_W_N_245_INT\ : std_logic;
signal \U_MD7AndNet\ : std_logic;
signal \U_MD7LegalizeSB_DFFNet\ : std_logic;
signal \U_ROMEN1_NLegalizeSB_DFFNet\ : std_logic;
signal \ROMEN2_N_c\ : std_logic;
signal \CASEN_N_padLegalizeSB_DFFNet\ : std_logic;
signal \CXXXOUT_padLegalizeSB_DFFNet\ : std_logic;
signal \EN80_N_padLegalizeSB_DFFNet\ : std_logic;
signal \ROMEN2_N_padLegalizeSB_DFFNet\ : std_logic;
signal \FXXX_N_N_8\ : std_logic;
signal \D_FXXX_cascade_\ : std_logic;
signal \D2_6_N_148\ : std_logic;
signal \C8_FXX_cascade_\ : std_logic;
signal \INTC8ACC\ : std_logic;
signal \CXXX_cascade_\ : std_logic;
signal n966 : std_logic;
signal \CXXX\ : std_logic;
signal \U_MMU_ROMEN.n7\ : std_logic;
signal \U_MMU_ROMEN.n4\ : std_logic;
signal \ROMEN1_N_INT\ : std_logic;
signal \INH_N_c\ : std_logic;
signal \CXXXOUT_c\ : std_logic;
signal \U_ADDR_DECODER.n2654\ : std_logic;
signal \EN80_N_c\ : std_logic;
signal n907 : std_logic;
signal \CASEN_N_c\ : std_logic;
signal \HIRES\ : std_logic;
signal \U_MMU_SELMB.n2572\ : std_logic;
signal \U_MMU_SELMB.n2610\ : std_logic;
signal \HIRES_cascade_\ : std_logic;
signal \WRPROT\ : std_logic;
signal \U_MMU_SOFT_SWITCHES_C08X.OUT_FST_ACC\ : std_logic;
signal \U_MMU_SOFT_SWITCHES_C08X.OUT_WREN\ : std_logic;
signal \INVU_MMU_SOFT_SWITCHES_C08X.OUT_FST_ACC_27C_net\ : std_logic;
signal \U_MMU_SELMB.n2516\ : std_logic;
signal \PG2\ : std_logic;
signal \SELMB_N\ : std_logic;
signal \D_PHI_0\ : std_logic;
signal \UMMU_INTERNALS.n1605_cascade_\ : std_logic;
signal \INTC8EN\ : std_logic;
signal \U_MMU_HOLD_TIME.SHIFT_REGISTER_1\ : std_logic;
signal \U_MMU_HOLD_TIME.SHIFT_REGISTER_0\ : std_logic;
signal n2596 : std_logic;
signal n911 : std_logic;
signal \RDRAM\ : std_logic;
signal \U_MMU_MD7.n2658_cascade_\ : std_logic;
signal \U_MMU_MD7.n2\ : std_logic;
signal \U_MMU_MD7.n2710\ : std_logic;
signal \UNGATED_MD7\ : std_logic;
signal \U_MMU_MD7.n2707\ : std_logic;
signal \BANK2\ : std_logic;
signal \INVU_MMU_SOFT_SWITCHES_C08X.BANK2_30C_net\ : std_logic;
signal \RDROM\ : std_logic;
signal \INVU_MMU_SOFT_SWITCHES_C08X.RDROM_31C_net\ : std_logic;
signal \INTC300_N_cascade_\ : std_logic;
signal \INTC3ACC_N_N_175\ : std_logic;
signal \U_MMU_RA.MMU_RA_MUX.D_Q3\ : std_logic;
signal \U_MMU_RA.MMU_RA_MUX.U_DRAM_HOLD_TIME.Q3_SHIFT_REGISTER_0\ : std_logic;
signal \U_MMU_RA.MMU_RA_MUX.U_DRAM_HOLD_TIME.Q3_SHIFT_REGISTER_1\ : std_logic;
signal n2584 : std_logic;
signal \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.n937\ : std_logic;
signal \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.n2532\ : std_logic;
signal \ALTSTKZP_cascade_\ : std_logic;
signal \INTC300_N\ : std_logic;
signal \U_MMU_MD7.n5\ : std_logic;
signal \FLG1\ : std_logic;
signal \ALTSTKZP\ : std_logic;
signal \SELMB_N_N_137_cascade_\ : std_logic;
signal \D_FXXX\ : std_logic;
signal \U_MMU_SELMB.SELMB_N_N_136\ : std_logic;
signal \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.n938\ : std_logic;
signal \DXXX_N_N_13\ : std_logic;
signal \BANK1\ : std_logic;
signal \ORA_pad_6AndNet\ : std_logic;
signal \ORA_pad_7AndNet\ : std_logic;
signal \KBD_N_padLegalizeSB_DFFNet\ : std_logic;
signal \ORA_pad_6LegalizeSB_DFFNet\ : std_logic;
signal \ORA_pad_7LegalizeSB_DFFNet\ : std_logic;
signal \CENROM1\ : std_logic;
signal \PENIO_N\ : std_logic;
signal \PENIO_N_cascade_\ : std_logic;
signal \U_MMU_MD7.n4\ : std_logic;
signal \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.n2570_cascade_\ : std_logic;
signal \EN80VID\ : std_logic;
signal n927 : std_logic;
signal \C8_FXX\ : std_logic;
signal \n927_cascade_\ : std_logic;
signal \UMMU_INTERNALS.n2616_cascade_\ : std_logic;
signal \UMMU_INTERNALS.n2622\ : std_logic;
signal \UNGATED_RA_6\ : std_logic;
signal \KBD_N_c\ : std_logic;
signal \UNGATED_RA_7\ : std_logic;
signal \U_MMU_RA.MMU_RA_MUX.U_DRAM_HOLD_TIME.PRAS_N_SHIFT_REGISTER_0\ : std_logic;
signal \U_MMU_RA.MMU_RA_MUX.U_DRAM_HOLD_TIME.PRAS_N_SHIFT_REGISTER_1\ : std_logic;
signal \A_c_14\ : std_logic;
signal \A_c_15\ : std_logic;
signal \U_MMU_MPON.n2521\ : std_logic;
signal \U_MMU_MPON.n2602_cascade_\ : std_logic;
signal \U_ADDR_DECODER.MC0XX_N_N_20\ : std_logic;
signal \MC0XX_N_cascade_\ : std_logic;
signal n2576 : std_logic;
signal \n1226_cascade_\ : std_logic;
signal \LATCHED_MC05X_N\ : std_logic;
signal n933 : std_logic;
signal \UMMU_INTERNALS.n2580\ : std_logic;
signal n2520 : std_logic;
signal \MA12_N_209\ : std_logic;
signal \U_MMU_RA.MMU_RA_MUX.COMBINED_RAS_N_cascade_\ : std_logic;
signal \A_c_12\ : std_logic;
signal \UNGATED_RA_4\ : std_logic;
signal \U_MMU_RA.MMU_RA_MUX.U_DRAM_HOLD_TIME.PRAS_N_SHIFT_REGISTER_2\ : std_logic;
signal \DELAY_CLK\ : std_logic;
signal \U_ADDR_DECODER.S_0XXX_N\ : std_logic;
signal \n953_cascade_\ : std_logic;
signal \DEV0_N\ : std_logic;
signal n953 : std_logic;
signal \ENABLE_N_cascade_\ : std_logic;
signal n912 : std_logic;
signal \MC0XX_N\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U_ADDR_DECODER.n44\ : std_logic;
signal \MD7_ENABLE_N_N_6\ : std_logic;
signal \A_c_13\ : std_logic;
signal \A_c_5\ : std_logic;
signal \UNGATED_RA_5\ : std_logic;
signal \A_c_4\ : std_logic;
signal \U_ADDR_DECODER.n9\ : std_logic;
signal \U_MMU_MPON.n13\ : std_logic;
signal \A_c_8\ : std_logic;
signal n626 : std_logic;
signal \U_MMU_MPON.M5_2\ : std_logic;
signal \U_MMU_MPON.M5_7\ : std_logic;
signal \U_MMU_MPON.DELTA_01XX_N\ : std_logic;
signal n2523 : std_logic;
signal \R_W_N_c\ : std_logic;
signal \n2523_cascade_\ : std_logic;
signal \U_ADDR_DECODER.n7\ : std_logic;
signal n906 : std_logic;
signal \INVU_MMU_RA.MMU_RA_MUX.RA_ENABLE_N_22C_net\ : std_logic;
signal \U_MMU_RA.MMU_RA_MUX.RA_ENABLE_N_N_215\ : std_logic;
signal \RA_ENABLE_N\ : std_logic;
signal \ORA_pad_3AndNet\ : std_logic;
signal \ORA_pad_4AndNet\ : std_logic;
signal \ORA_pad_5AndNet\ : std_logic;
signal \ORA_pad_3LegalizeSB_DFFNet\ : std_logic;
signal \ORA_pad_4LegalizeSB_DFFNet\ : std_logic;
signal \ORA_pad_5LegalizeSB_DFFNet\ : std_logic;
signal \Q3_c\ : std_logic;
signal \PHI_0_c\ : std_logic;
signal n2620 : std_logic;
signal n949 : std_logic;
signal \n15_cascade_\ : std_logic;
signal n16 : std_logic;
signal \ENABLE_N\ : std_logic;
signal \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.n2566\ : std_logic;
signal \MPON_N\ : std_logic;
signal \FLG2\ : std_logic;
signal \A_c_11\ : std_logic;
signal \A_c_3\ : std_logic;
signal \UNGATED_RA_3\ : std_logic;
signal \A_c_9\ : std_logic;
signal \A_c_0\ : std_logic;
signal \UNGATED_RA_0\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_1\ : std_logic;
signal \UNGATED_RA_1\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U_MMU_RA.MMU_RA_MUX.D_RAS_N\ : std_logic;
signal \PRAS_N_c\ : std_logic;
signal \A_c_10\ : std_logic;
signal \UNGATED_RA_2\ : std_logic;
signal \ORA_pad_0AndNet\ : std_logic;
signal \ORA_pad_1AndNet\ : std_logic;
signal \RA_ENABLE_N_N_2\ : std_logic;
signal \ORA_pad_2AndNet\ : std_logic;
signal \ORA_pad_0LegalizeSB_DFFNet\ : std_logic;
signal \ORA_pad_1LegalizeSB_DFFNet\ : std_logic;
signal \ORA_pad_2LegalizeSB_DFFNet\ : std_logic;
signal \internalOscilatorOutputNet\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \PHI_0_wire\ : std_logic;
signal \ORA_wire\ : std_logic_vector(7 downto 0);
signal \Q3_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(15 downto 0);
signal \CXXXOUT_wire\ : std_logic;
signal \DMA_N_wire\ : std_logic;
signal \KBD_N_wire\ : std_logic;
signal \EN80_N_wire\ : std_logic;
signal \R_W_N_wire\ : std_logic;
signal \CASEN_N_wire\ : std_logic;
signal \INH_N_wire\ : std_logic;
signal \ROMEN2_N_wire\ : std_logic;
signal \PRAS_N_wire\ : std_logic;

begin
    \PHI_0_wire\ <= PHI_0;
    ORA <= \ORA_wire\;
    \Q3_wire\ <= Q3;
    \A_wire\ <= A;
    CXXXOUT <= \CXXXOUT_wire\;
    \DMA_N_wire\ <= DMA_N;
    KBD_N <= \KBD_N_wire\;
    EN80_N <= \EN80_N_wire\;
    \R_W_N_wire\ <= R_W_N;
    CASEN_N <= \CASEN_N_wire\;
    \INH_N_wire\ <= INH_N;
    ROMEN2_N <= \ROMEN2_N_wire\;
    \PRAS_N_wire\ <= PRAS_N;

    \PHI_0_pad_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__6165\,
            GLOBALBUFFEROUTPUT => \PHI_0_c\
        );

    \PHI_0_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6167\,
            DIN => \N__6166\,
            DOUT => \N__6165\,
            PACKAGEPIN => \PHI_0_wire\
        );

    \PHI_0_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6167\,
            PADOUT => \N__6166\,
            PADIN => \N__6165\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ORA_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6156\,
            DIN => \N__6155\,
            DOUT => \N__6154\,
            PACKAGEPIN => \ORA_wire\(7)
        );

    \ORA_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6156\,
            PADOUT => \N__6155\,
            PADIN => \N__6154\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2915\,
            DIN0 => OPEN,
            DOUT0 => \N__3266\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Q3_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6147\,
            DIN => \N__6146\,
            DOUT => \N__6145\,
            PACKAGEPIN => \Q3_wire\
        );

    \Q3_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6147\,
            PADOUT => \N__6146\,
            PADIN => \N__6145\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \Q3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6138\,
            DIN => \N__6137\,
            DOUT => \N__6136\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6138\,
            PADOUT => \N__6137\,
            PADIN => \N__6136\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CXXXOUT_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6129\,
            DIN => \N__6128\,
            DOUT => \N__6127\,
            PACKAGEPIN => \CXXXOUT_wire\
        );

    \CXXXOUT_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6129\,
            PADOUT => \N__6128\,
            PADIN => \N__6127\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2216\,
            DIN0 => OPEN,
            DOUT0 => \N__2396\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_N_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6120\,
            DIN => \N__6119\,
            DOUT => \N__6118\,
            PACKAGEPIN => \DMA_N_wire\
        );

    \DMA_N_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6120\,
            PADOUT => \N__6119\,
            PADIN => \N__6118\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DMA_N_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \KBD_N_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6111\,
            DIN => \N__6110\,
            DOUT => \N__6109\,
            PACKAGEPIN => \KBD_N_wire\
        );

    \KBD_N_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6111\,
            PADOUT => \N__6110\,
            PADIN => \N__6109\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2909\,
            DIN0 => OPEN,
            DOUT0 => \N__2984\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_pad_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6102\,
            DIN => \N__6101\,
            DOUT => \N__6100\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_pad_13_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6102\,
            PADOUT => \N__6101\,
            PADIN => \N__6100\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \EN80_N_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6093\,
            DIN => \N__6092\,
            DOUT => \N__6091\,
            PACKAGEPIN => \EN80_N_wire\
        );

    \EN80_N_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6093\,
            PADOUT => \N__6092\,
            PADIN => \N__6091\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2210\,
            DIN0 => OPEN,
            DOUT0 => \N__2369\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ORA_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6084\,
            DIN => \N__6083\,
            DOUT => \N__6082\,
            PACKAGEPIN => \ORA_wire\(4)
        );

    \ORA_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6084\,
            PADOUT => \N__6083\,
            PADIN => \N__6082\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4322\,
            DIN0 => OPEN,
            DOUT0 => \N__3323\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6075\,
            DIN => \N__6074\,
            DOUT => \N__6073\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6075\,
            PADOUT => \N__6074\,
            PADIN => \N__6073\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ORA_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6066\,
            DIN => \N__6065\,
            DOUT => \N__6064\,
            PACKAGEPIN => \ORA_wire\(0)
        );

    \ORA_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6066\,
            PADOUT => \N__6065\,
            PADIN => \N__6064\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4358\,
            DIN0 => OPEN,
            DOUT0 => \N__5012\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ORA_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6057\,
            DIN => \N__6056\,
            DOUT => \N__6055\,
            PACKAGEPIN => \ORA_wire\(5)
        );

    \ORA_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6057\,
            PADOUT => \N__6056\,
            PADIN => \N__6055\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4316\,
            DIN0 => OPEN,
            DOUT0 => \N__3545\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \R_W_N_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6048\,
            DIN => \N__6047\,
            DOUT => \N__6046\,
            PACKAGEPIN => \R_W_N_wire\
        );

    \R_W_N_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6048\,
            PADOUT => \N__6047\,
            PADIN => \N__6046\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \R_W_N_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6039\,
            DIN => \N__6038\,
            DOUT => \N__6037\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6039\,
            PADOUT => \N__6038\,
            PADIN => \N__6037\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_pad_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6030\,
            DIN => \N__6029\,
            DOUT => \N__6028\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_pad_10_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6030\,
            PADOUT => \N__6029\,
            PADIN => \N__6028\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ORA_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6021\,
            DIN => \N__6020\,
            DOUT => \N__6019\,
            PACKAGEPIN => \ORA_wire\(1)
        );

    \ORA_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6021\,
            PADOUT => \N__6020\,
            PADIN => \N__6019\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5840\,
            DIN0 => OPEN,
            DOUT0 => \N__4772\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6012\,
            DIN => \N__6011\,
            DOUT => \N__6010\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6012\,
            PADOUT => \N__6011\,
            PADIN => \N__6010\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_pad_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6003\,
            DIN => \N__6002\,
            DOUT => \N__6001\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_pad_14_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__6003\,
            PADOUT => \N__6002\,
            PADIN => \N__6001\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ORA_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5994\,
            DIN => \N__5993\,
            DOUT => \N__5992\,
            PACKAGEPIN => \ORA_wire\(6)
        );

    \ORA_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5994\,
            PADOUT => \N__5993\,
            PADIN => \N__5992\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2921\,
            DIN0 => OPEN,
            DOUT0 => \N__2996\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5985\,
            DIN => \N__5984\,
            DOUT => \N__5983\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5985\,
            PADOUT => \N__5984\,
            PADIN => \N__5983\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_pad_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5976\,
            DIN => \N__5975\,
            DOUT => \N__5974\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_pad_9_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5976\,
            PADOUT => \N__5975\,
            PADIN => \N__5974\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_pad_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5967\,
            DIN => \N__5966\,
            DOUT => \N__5965\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_pad_11_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5967\,
            PADOUT => \N__5966\,
            PADIN => \N__5965\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ORA_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5958\,
            DIN => \N__5957\,
            DOUT => \N__5956\,
            PACKAGEPIN => \ORA_wire\(2)
        );

    \ORA_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5958\,
            PADOUT => \N__5957\,
            PADIN => \N__5956\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5786\,
            DIN0 => OPEN,
            DOUT0 => \N__4370\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5949\,
            DIN => \N__5948\,
            DOUT => \N__5947\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5949\,
            PADOUT => \N__5948\,
            PADIN => \N__5947\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_pad_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5940\,
            DIN => \N__5939\,
            DOUT => \N__5938\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_pad_15_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5940\,
            PADOUT => \N__5939\,
            PADIN => \N__5938\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_pad_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5931\,
            DIN => \N__5930\,
            DOUT => \N__5929\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_pad_8_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5931\,
            PADOUT => \N__5930\,
            PADIN => \N__5929\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASEN_N_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5922\,
            DIN => \N__5921\,
            DOUT => \N__5920\,
            PACKAGEPIN => \CASEN_N_wire\
        );

    \CASEN_N_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5922\,
            PADOUT => \N__5921\,
            PADIN => \N__5920\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2222\,
            DIN0 => OPEN,
            DOUT0 => \N__2342\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_pad_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5913\,
            DIN => \N__5912\,
            DOUT => \N__5911\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_pad_12_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5913\,
            PADOUT => \N__5912\,
            PADIN => \N__5911\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ORA_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5904\,
            DIN => \N__5903\,
            DOUT => \N__5902\,
            PACKAGEPIN => \ORA_wire\(3)
        );

    \ORA_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5904\,
            PADOUT => \N__5903\,
            PADIN => \N__5902\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4328\,
            DIN0 => OPEN,
            DOUT0 => \N__5252\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5895\,
            DIN => \N__5894\,
            DOUT => \N__5893\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5895\,
            PADOUT => \N__5894\,
            PADIN => \N__5893\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \INH_N_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5886\,
            DIN => \N__5885\,
            DOUT => \N__5884\,
            PACKAGEPIN => \INH_N_wire\
        );

    \INH_N_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5886\,
            PADOUT => \N__5885\,
            PADIN => \N__5884\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \INH_N_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ROMEN2_N_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5877\,
            DIN => \N__5876\,
            DOUT => \N__5875\,
            PACKAGEPIN => \ROMEN2_N_wire\
        );

    \ROMEN2_N_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5877\,
            PADOUT => \N__5876\,
            PADIN => \N__5875\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2204\,
            DIN0 => OPEN,
            DOUT0 => \N__2234\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5868\,
            DIN => \N__5867\,
            DOUT => \N__5866\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5868\,
            PADOUT => \N__5867\,
            PADIN => \N__5866\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PRAS_N_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5859\,
            DIN => \N__5858\,
            DOUT => \N__5857\,
            PACKAGEPIN => \PRAS_N_wire\
        );

    \PRAS_N_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__5859\,
            PADOUT => \N__5858\,
            PADIN => \N__5857\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \PRAS_N_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1408\ : IoInMux
    port map (
            O => \N__5840\,
            I => \N__5837\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__5837\,
            I => \ORA_pad_1AndNet\
        );

    \I__1406\ : InMux
    port map (
            O => \N__5834\,
            I => \N__5825\
        );

    \I__1405\ : InMux
    port map (
            O => \N__5833\,
            I => \N__5825\
        );

    \I__1404\ : InMux
    port map (
            O => \N__5832\,
            I => \N__5818\
        );

    \I__1403\ : InMux
    port map (
            O => \N__5831\,
            I => \N__5818\
        );

    \I__1402\ : InMux
    port map (
            O => \N__5830\,
            I => \N__5818\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__5825\,
            I => \N__5812\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__5818\,
            I => \N__5809\
        );

    \I__1399\ : InMux
    port map (
            O => \N__5817\,
            I => \N__5802\
        );

    \I__1398\ : InMux
    port map (
            O => \N__5816\,
            I => \N__5802\
        );

    \I__1397\ : InMux
    port map (
            O => \N__5815\,
            I => \N__5802\
        );

    \I__1396\ : Span4Mux_v
    port map (
            O => \N__5812\,
            I => \N__5799\
        );

    \I__1395\ : Span4Mux_v
    port map (
            O => \N__5809\,
            I => \N__5796\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__5802\,
            I => \N__5793\
        );

    \I__1393\ : Odrv4
    port map (
            O => \N__5799\,
            I => \RA_ENABLE_N_N_2\
        );

    \I__1392\ : Odrv4
    port map (
            O => \N__5796\,
            I => \RA_ENABLE_N_N_2\
        );

    \I__1391\ : Odrv12
    port map (
            O => \N__5793\,
            I => \RA_ENABLE_N_N_2\
        );

    \I__1390\ : IoInMux
    port map (
            O => \N__5786\,
            I => \N__5783\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__5783\,
            I => \ORA_pad_2AndNet\
        );

    \I__1388\ : InMux
    port map (
            O => \N__5780\,
            I => \N__5777\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__5777\,
            I => \ORA_pad_0LegalizeSB_DFFNet\
        );

    \I__1386\ : InMux
    port map (
            O => \N__5774\,
            I => \N__5771\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__5771\,
            I => \ORA_pad_1LegalizeSB_DFFNet\
        );

    \I__1384\ : InMux
    port map (
            O => \N__5768\,
            I => \N__5765\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__5765\,
            I => \ORA_pad_2LegalizeSB_DFFNet\
        );

    \I__1382\ : ClkMux
    port map (
            O => \N__5762\,
            I => \N__5759\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__5759\,
            I => \N__5755\
        );

    \I__1380\ : ClkMux
    port map (
            O => \N__5758\,
            I => \N__5752\
        );

    \I__1379\ : Span4Mux_h
    port map (
            O => \N__5755\,
            I => \N__5746\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__5752\,
            I => \N__5746\
        );

    \I__1377\ : ClkMux
    port map (
            O => \N__5751\,
            I => \N__5743\
        );

    \I__1376\ : Span4Mux_h
    port map (
            O => \N__5746\,
            I => \N__5736\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__5743\,
            I => \N__5736\
        );

    \I__1374\ : ClkMux
    port map (
            O => \N__5742\,
            I => \N__5733\
        );

    \I__1373\ : ClkMux
    port map (
            O => \N__5741\,
            I => \N__5729\
        );

    \I__1372\ : Span4Mux_h
    port map (
            O => \N__5736\,
            I => \N__5724\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__5733\,
            I => \N__5724\
        );

    \I__1370\ : ClkMux
    port map (
            O => \N__5732\,
            I => \N__5721\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__5729\,
            I => \N__5718\
        );

    \I__1368\ : Span4Mux_h
    port map (
            O => \N__5724\,
            I => \N__5713\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__5721\,
            I => \N__5713\
        );

    \I__1366\ : Span12Mux_h
    port map (
            O => \N__5718\,
            I => \N__5710\
        );

    \I__1365\ : Sp12to4
    port map (
            O => \N__5713\,
            I => \N__5707\
        );

    \I__1364\ : Span12Mux_v
    port map (
            O => \N__5710\,
            I => \N__5704\
        );

    \I__1363\ : Span12Mux_h
    port map (
            O => \N__5707\,
            I => \N__5701\
        );

    \I__1362\ : Span12Mux_h
    port map (
            O => \N__5704\,
            I => \N__5696\
        );

    \I__1361\ : Span12Mux_v
    port map (
            O => \N__5701\,
            I => \N__5696\
        );

    \I__1360\ : Odrv12
    port map (
            O => \N__5696\,
            I => \internalOscilatorOutputNet\
        );

    \I__1359\ : InMux
    port map (
            O => \N__5693\,
            I => \N__5690\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__5690\,
            I => \N__5687\
        );

    \I__1357\ : Odrv12
    port map (
            O => \N__5687\,
            I => n2620
        );

    \I__1356\ : InMux
    port map (
            O => \N__5684\,
            I => \N__5681\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__5681\,
            I => n949
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__5678\,
            I => \n15_cascade_\
        );

    \I__1353\ : InMux
    port map (
            O => \N__5675\,
            I => \N__5672\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__5672\,
            I => \N__5669\
        );

    \I__1351\ : Odrv4
    port map (
            O => \N__5669\,
            I => n16
        );

    \I__1350\ : InMux
    port map (
            O => \N__5666\,
            I => \N__5660\
        );

    \I__1349\ : InMux
    port map (
            O => \N__5665\,
            I => \N__5657\
        );

    \I__1348\ : InMux
    port map (
            O => \N__5664\,
            I => \N__5654\
        );

    \I__1347\ : InMux
    port map (
            O => \N__5663\,
            I => \N__5651\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__5660\,
            I => \N__5647\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__5657\,
            I => \N__5644\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__5654\,
            I => \N__5641\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__5651\,
            I => \N__5638\
        );

    \I__1342\ : InMux
    port map (
            O => \N__5650\,
            I => \N__5635\
        );

    \I__1341\ : Span4Mux_v
    port map (
            O => \N__5647\,
            I => \N__5630\
        );

    \I__1340\ : Span4Mux_v
    port map (
            O => \N__5644\,
            I => \N__5630\
        );

    \I__1339\ : Span4Mux_v
    port map (
            O => \N__5641\,
            I => \N__5623\
        );

    \I__1338\ : Span4Mux_v
    port map (
            O => \N__5638\,
            I => \N__5623\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__5635\,
            I => \N__5623\
        );

    \I__1336\ : Odrv4
    port map (
            O => \N__5630\,
            I => \ENABLE_N\
        );

    \I__1335\ : Odrv4
    port map (
            O => \N__5623\,
            I => \ENABLE_N\
        );

    \I__1334\ : InMux
    port map (
            O => \N__5618\,
            I => \N__5615\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__5615\,
            I => \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.n2566\
        );

    \I__1332\ : CascadeMux
    port map (
            O => \N__5612\,
            I => \N__5608\
        );

    \I__1331\ : SRMux
    port map (
            O => \N__5611\,
            I => \N__5603\
        );

    \I__1330\ : InMux
    port map (
            O => \N__5608\,
            I => \N__5600\
        );

    \I__1329\ : CascadeMux
    port map (
            O => \N__5607\,
            I => \N__5596\
        );

    \I__1328\ : CascadeMux
    port map (
            O => \N__5606\,
            I => \N__5587\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__5603\,
            I => \N__5584\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__5600\,
            I => \N__5581\
        );

    \I__1325\ : InMux
    port map (
            O => \N__5599\,
            I => \N__5578\
        );

    \I__1324\ : InMux
    port map (
            O => \N__5596\,
            I => \N__5575\
        );

    \I__1323\ : InMux
    port map (
            O => \N__5595\,
            I => \N__5572\
        );

    \I__1322\ : SRMux
    port map (
            O => \N__5594\,
            I => \N__5569\
        );

    \I__1321\ : SRMux
    port map (
            O => \N__5593\,
            I => \N__5566\
        );

    \I__1320\ : InMux
    port map (
            O => \N__5592\,
            I => \N__5563\
        );

    \I__1319\ : InMux
    port map (
            O => \N__5591\,
            I => \N__5560\
        );

    \I__1318\ : InMux
    port map (
            O => \N__5590\,
            I => \N__5557\
        );

    \I__1317\ : InMux
    port map (
            O => \N__5587\,
            I => \N__5554\
        );

    \I__1316\ : Span4Mux_v
    port map (
            O => \N__5584\,
            I => \N__5551\
        );

    \I__1315\ : Span4Mux_h
    port map (
            O => \N__5581\,
            I => \N__5538\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__5578\,
            I => \N__5538\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__5575\,
            I => \N__5538\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__5572\,
            I => \N__5538\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__5569\,
            I => \N__5538\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__5566\,
            I => \N__5538\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__5563\,
            I => \N__5528\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__5560\,
            I => \N__5528\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__5557\,
            I => \N__5528\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__5554\,
            I => \N__5528\
        );

    \I__1305\ : Span4Mux_h
    port map (
            O => \N__5551\,
            I => \N__5522\
        );

    \I__1304\ : Span4Mux_v
    port map (
            O => \N__5538\,
            I => \N__5522\
        );

    \I__1303\ : InMux
    port map (
            O => \N__5537\,
            I => \N__5519\
        );

    \I__1302\ : Span4Mux_v
    port map (
            O => \N__5528\,
            I => \N__5516\
        );

    \I__1301\ : InMux
    port map (
            O => \N__5527\,
            I => \N__5513\
        );

    \I__1300\ : Span4Mux_h
    port map (
            O => \N__5522\,
            I => \N__5510\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__5519\,
            I => \N__5507\
        );

    \I__1298\ : Span4Mux_h
    port map (
            O => \N__5516\,
            I => \N__5502\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__5513\,
            I => \N__5502\
        );

    \I__1296\ : Odrv4
    port map (
            O => \N__5510\,
            I => \MPON_N\
        );

    \I__1295\ : Odrv12
    port map (
            O => \N__5507\,
            I => \MPON_N\
        );

    \I__1294\ : Odrv4
    port map (
            O => \N__5502\,
            I => \MPON_N\
        );

    \I__1293\ : InMux
    port map (
            O => \N__5495\,
            I => \N__5492\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__5492\,
            I => \N__5489\
        );

    \I__1291\ : Span4Mux_v
    port map (
            O => \N__5489\,
            I => \N__5484\
        );

    \I__1290\ : InMux
    port map (
            O => \N__5488\,
            I => \N__5481\
        );

    \I__1289\ : CascadeMux
    port map (
            O => \N__5487\,
            I => \N__5478\
        );

    \I__1288\ : Sp12to4
    port map (
            O => \N__5484\,
            I => \N__5473\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__5481\,
            I => \N__5473\
        );

    \I__1286\ : InMux
    port map (
            O => \N__5478\,
            I => \N__5470\
        );

    \I__1285\ : Odrv12
    port map (
            O => \N__5473\,
            I => \FLG2\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__5470\,
            I => \FLG2\
        );

    \I__1283\ : InMux
    port map (
            O => \N__5465\,
            I => \N__5460\
        );

    \I__1282\ : CascadeMux
    port map (
            O => \N__5464\,
            I => \N__5456\
        );

    \I__1281\ : InMux
    port map (
            O => \N__5463\,
            I => \N__5453\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__5460\,
            I => \N__5450\
        );

    \I__1279\ : InMux
    port map (
            O => \N__5459\,
            I => \N__5446\
        );

    \I__1278\ : InMux
    port map (
            O => \N__5456\,
            I => \N__5443\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__5453\,
            I => \N__5439\
        );

    \I__1276\ : Span4Mux_v
    port map (
            O => \N__5450\,
            I => \N__5436\
        );

    \I__1275\ : InMux
    port map (
            O => \N__5449\,
            I => \N__5433\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__5446\,
            I => \N__5430\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__5443\,
            I => \N__5427\
        );

    \I__1272\ : InMux
    port map (
            O => \N__5442\,
            I => \N__5424\
        );

    \I__1271\ : Span4Mux_h
    port map (
            O => \N__5439\,
            I => \N__5421\
        );

    \I__1270\ : Span4Mux_h
    port map (
            O => \N__5436\,
            I => \N__5416\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__5433\,
            I => \N__5416\
        );

    \I__1268\ : Span12Mux_h
    port map (
            O => \N__5430\,
            I => \N__5413\
        );

    \I__1267\ : Span12Mux_h
    port map (
            O => \N__5427\,
            I => \N__5408\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__5424\,
            I => \N__5408\
        );

    \I__1265\ : Span4Mux_v
    port map (
            O => \N__5421\,
            I => \N__5405\
        );

    \I__1264\ : Span4Mux_h
    port map (
            O => \N__5416\,
            I => \N__5402\
        );

    \I__1263\ : Odrv12
    port map (
            O => \N__5413\,
            I => \A_c_11\
        );

    \I__1262\ : Odrv12
    port map (
            O => \N__5408\,
            I => \A_c_11\
        );

    \I__1261\ : Odrv4
    port map (
            O => \N__5405\,
            I => \A_c_11\
        );

    \I__1260\ : Odrv4
    port map (
            O => \N__5402\,
            I => \A_c_11\
        );

    \I__1259\ : InMux
    port map (
            O => \N__5393\,
            I => \N__5387\
        );

    \I__1258\ : InMux
    port map (
            O => \N__5392\,
            I => \N__5382\
        );

    \I__1257\ : InMux
    port map (
            O => \N__5391\,
            I => \N__5382\
        );

    \I__1256\ : CascadeMux
    port map (
            O => \N__5390\,
            I => \N__5379\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__5387\,
            I => \N__5371\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__5382\,
            I => \N__5371\
        );

    \I__1253\ : InMux
    port map (
            O => \N__5379\,
            I => \N__5366\
        );

    \I__1252\ : InMux
    port map (
            O => \N__5378\,
            I => \N__5366\
        );

    \I__1251\ : InMux
    port map (
            O => \N__5377\,
            I => \N__5360\
        );

    \I__1250\ : InMux
    port map (
            O => \N__5376\,
            I => \N__5357\
        );

    \I__1249\ : Span4Mux_v
    port map (
            O => \N__5371\,
            I => \N__5349\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__5366\,
            I => \N__5349\
        );

    \I__1247\ : InMux
    port map (
            O => \N__5365\,
            I => \N__5346\
        );

    \I__1246\ : InMux
    port map (
            O => \N__5364\,
            I => \N__5343\
        );

    \I__1245\ : CascadeMux
    port map (
            O => \N__5363\,
            I => \N__5340\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__5360\,
            I => \N__5334\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__5357\,
            I => \N__5334\
        );

    \I__1242\ : InMux
    port map (
            O => \N__5356\,
            I => \N__5331\
        );

    \I__1241\ : InMux
    port map (
            O => \N__5355\,
            I => \N__5328\
        );

    \I__1240\ : InMux
    port map (
            O => \N__5354\,
            I => \N__5325\
        );

    \I__1239\ : Span4Mux_v
    port map (
            O => \N__5349\,
            I => \N__5322\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__5346\,
            I => \N__5317\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__5343\,
            I => \N__5317\
        );

    \I__1236\ : InMux
    port map (
            O => \N__5340\,
            I => \N__5314\
        );

    \I__1235\ : InMux
    port map (
            O => \N__5339\,
            I => \N__5310\
        );

    \I__1234\ : Span4Mux_v
    port map (
            O => \N__5334\,
            I => \N__5306\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__5331\,
            I => \N__5301\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__5328\,
            I => \N__5301\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__5325\,
            I => \N__5298\
        );

    \I__1230\ : Span4Mux_h
    port map (
            O => \N__5322\,
            I => \N__5291\
        );

    \I__1229\ : Span4Mux_v
    port map (
            O => \N__5317\,
            I => \N__5291\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__5314\,
            I => \N__5291\
        );

    \I__1227\ : CascadeMux
    port map (
            O => \N__5313\,
            I => \N__5288\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__5310\,
            I => \N__5285\
        );

    \I__1225\ : InMux
    port map (
            O => \N__5309\,
            I => \N__5282\
        );

    \I__1224\ : Span4Mux_h
    port map (
            O => \N__5306\,
            I => \N__5275\
        );

    \I__1223\ : Span4Mux_v
    port map (
            O => \N__5301\,
            I => \N__5275\
        );

    \I__1222\ : Span4Mux_v
    port map (
            O => \N__5298\,
            I => \N__5275\
        );

    \I__1221\ : Span4Mux_v
    port map (
            O => \N__5291\,
            I => \N__5272\
        );

    \I__1220\ : InMux
    port map (
            O => \N__5288\,
            I => \N__5269\
        );

    \I__1219\ : Span12Mux_v
    port map (
            O => \N__5285\,
            I => \N__5258\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__5282\,
            I => \N__5258\
        );

    \I__1217\ : Sp12to4
    port map (
            O => \N__5275\,
            I => \N__5258\
        );

    \I__1216\ : Sp12to4
    port map (
            O => \N__5272\,
            I => \N__5258\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__5269\,
            I => \N__5258\
        );

    \I__1214\ : Span12Mux_h
    port map (
            O => \N__5258\,
            I => \N__5255\
        );

    \I__1213\ : Odrv12
    port map (
            O => \N__5255\,
            I => \A_c_3\
        );

    \I__1212\ : IoInMux
    port map (
            O => \N__5252\,
            I => \N__5249\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__5249\,
            I => \N__5246\
        );

    \I__1210\ : Sp12to4
    port map (
            O => \N__5246\,
            I => \N__5243\
        );

    \I__1209\ : Odrv12
    port map (
            O => \N__5243\,
            I => \UNGATED_RA_3\
        );

    \I__1208\ : CascadeMux
    port map (
            O => \N__5240\,
            I => \N__5236\
        );

    \I__1207\ : InMux
    port map (
            O => \N__5239\,
            I => \N__5233\
        );

    \I__1206\ : InMux
    port map (
            O => \N__5236\,
            I => \N__5228\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__5233\,
            I => \N__5225\
        );

    \I__1204\ : InMux
    port map (
            O => \N__5232\,
            I => \N__5222\
        );

    \I__1203\ : CascadeMux
    port map (
            O => \N__5231\,
            I => \N__5218\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__5228\,
            I => \N__5215\
        );

    \I__1201\ : Span4Mux_h
    port map (
            O => \N__5225\,
            I => \N__5210\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__5222\,
            I => \N__5210\
        );

    \I__1199\ : InMux
    port map (
            O => \N__5221\,
            I => \N__5207\
        );

    \I__1198\ : InMux
    port map (
            O => \N__5218\,
            I => \N__5204\
        );

    \I__1197\ : Span12Mux_s10_h
    port map (
            O => \N__5215\,
            I => \N__5201\
        );

    \I__1196\ : Span4Mux_v
    port map (
            O => \N__5210\,
            I => \N__5196\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__5207\,
            I => \N__5196\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__5204\,
            I => \N__5193\
        );

    \I__1193\ : Odrv12
    port map (
            O => \N__5201\,
            I => \A_c_9\
        );

    \I__1192\ : Odrv4
    port map (
            O => \N__5196\,
            I => \A_c_9\
        );

    \I__1191\ : Odrv12
    port map (
            O => \N__5193\,
            I => \A_c_9\
        );

    \I__1190\ : CascadeMux
    port map (
            O => \N__5186\,
            I => \N__5180\
        );

    \I__1189\ : InMux
    port map (
            O => \N__5185\,
            I => \N__5173\
        );

    \I__1188\ : CascadeMux
    port map (
            O => \N__5184\,
            I => \N__5163\
        );

    \I__1187\ : CascadeMux
    port map (
            O => \N__5183\,
            I => \N__5159\
        );

    \I__1186\ : InMux
    port map (
            O => \N__5180\,
            I => \N__5154\
        );

    \I__1185\ : InMux
    port map (
            O => \N__5179\,
            I => \N__5149\
        );

    \I__1184\ : InMux
    port map (
            O => \N__5178\,
            I => \N__5149\
        );

    \I__1183\ : InMux
    port map (
            O => \N__5177\,
            I => \N__5144\
        );

    \I__1182\ : InMux
    port map (
            O => \N__5176\,
            I => \N__5144\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__5173\,
            I => \N__5141\
        );

    \I__1180\ : InMux
    port map (
            O => \N__5172\,
            I => \N__5136\
        );

    \I__1179\ : InMux
    port map (
            O => \N__5171\,
            I => \N__5136\
        );

    \I__1178\ : InMux
    port map (
            O => \N__5170\,
            I => \N__5133\
        );

    \I__1177\ : InMux
    port map (
            O => \N__5169\,
            I => \N__5130\
        );

    \I__1176\ : InMux
    port map (
            O => \N__5168\,
            I => \N__5125\
        );

    \I__1175\ : InMux
    port map (
            O => \N__5167\,
            I => \N__5125\
        );

    \I__1174\ : InMux
    port map (
            O => \N__5166\,
            I => \N__5122\
        );

    \I__1173\ : InMux
    port map (
            O => \N__5163\,
            I => \N__5117\
        );

    \I__1172\ : InMux
    port map (
            O => \N__5162\,
            I => \N__5117\
        );

    \I__1171\ : InMux
    port map (
            O => \N__5159\,
            I => \N__5114\
        );

    \I__1170\ : InMux
    port map (
            O => \N__5158\,
            I => \N__5111\
        );

    \I__1169\ : InMux
    port map (
            O => \N__5157\,
            I => \N__5108\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__5154\,
            I => \N__5098\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__5149\,
            I => \N__5098\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__5144\,
            I => \N__5098\
        );

    \I__1165\ : Span4Mux_v
    port map (
            O => \N__5141\,
            I => \N__5093\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__5136\,
            I => \N__5093\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__5133\,
            I => \N__5082\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__5130\,
            I => \N__5082\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__5125\,
            I => \N__5082\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__5122\,
            I => \N__5082\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__5117\,
            I => \N__5082\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__5114\,
            I => \N__5077\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__5111\,
            I => \N__5077\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__5108\,
            I => \N__5074\
        );

    \I__1155\ : InMux
    port map (
            O => \N__5107\,
            I => \N__5071\
        );

    \I__1154\ : InMux
    port map (
            O => \N__5106\,
            I => \N__5068\
        );

    \I__1153\ : InMux
    port map (
            O => \N__5105\,
            I => \N__5064\
        );

    \I__1152\ : Span4Mux_v
    port map (
            O => \N__5098\,
            I => \N__5061\
        );

    \I__1151\ : Span4Mux_v
    port map (
            O => \N__5093\,
            I => \N__5058\
        );

    \I__1150\ : Span4Mux_v
    port map (
            O => \N__5082\,
            I => \N__5053\
        );

    \I__1149\ : Span4Mux_h
    port map (
            O => \N__5077\,
            I => \N__5053\
        );

    \I__1148\ : Span4Mux_v
    port map (
            O => \N__5074\,
            I => \N__5046\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__5071\,
            I => \N__5046\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__5068\,
            I => \N__5046\
        );

    \I__1145\ : InMux
    port map (
            O => \N__5067\,
            I => \N__5043\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__5064\,
            I => \N__5040\
        );

    \I__1143\ : Sp12to4
    port map (
            O => \N__5061\,
            I => \N__5035\
        );

    \I__1142\ : Sp12to4
    port map (
            O => \N__5058\,
            I => \N__5035\
        );

    \I__1141\ : Span4Mux_h
    port map (
            O => \N__5053\,
            I => \N__5028\
        );

    \I__1140\ : Span4Mux_v
    port map (
            O => \N__5046\,
            I => \N__5028\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__5043\,
            I => \N__5028\
        );

    \I__1138\ : Span12Mux_h
    port map (
            O => \N__5040\,
            I => \N__5025\
        );

    \I__1137\ : Span12Mux_h
    port map (
            O => \N__5035\,
            I => \N__5022\
        );

    \I__1136\ : Span4Mux_h
    port map (
            O => \N__5028\,
            I => \N__5019\
        );

    \I__1135\ : Odrv12
    port map (
            O => \N__5025\,
            I => \A_c_0\
        );

    \I__1134\ : Odrv12
    port map (
            O => \N__5022\,
            I => \A_c_0\
        );

    \I__1133\ : Odrv4
    port map (
            O => \N__5019\,
            I => \A_c_0\
        );

    \I__1132\ : IoInMux
    port map (
            O => \N__5012\,
            I => \N__5009\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__5009\,
            I => \N__5006\
        );

    \I__1130\ : Span12Mux_s11_v
    port map (
            O => \N__5006\,
            I => \N__5003\
        );

    \I__1129\ : Odrv12
    port map (
            O => \N__5003\,
            I => \UNGATED_RA_0\
        );

    \I__1128\ : InMux
    port map (
            O => \N__5000\,
            I => \N__4996\
        );

    \I__1127\ : InMux
    port map (
            O => \N__4999\,
            I => \N__4993\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__4996\,
            I => \N__4986\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__4993\,
            I => \N__4986\
        );

    \I__1124\ : InMux
    port map (
            O => \N__4992\,
            I => \N__4983\
        );

    \I__1123\ : InMux
    port map (
            O => \N__4991\,
            I => \N__4979\
        );

    \I__1122\ : Span4Mux_v
    port map (
            O => \N__4986\,
            I => \N__4974\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__4983\,
            I => \N__4974\
        );

    \I__1120\ : InMux
    port map (
            O => \N__4982\,
            I => \N__4971\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__4979\,
            I => \N__4967\
        );

    \I__1118\ : Span4Mux_v
    port map (
            O => \N__4974\,
            I => \N__4962\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__4971\,
            I => \N__4962\
        );

    \I__1116\ : CascadeMux
    port map (
            O => \N__4970\,
            I => \N__4959\
        );

    \I__1115\ : Span4Mux_h
    port map (
            O => \N__4967\,
            I => \N__4956\
        );

    \I__1114\ : Span4Mux_h
    port map (
            O => \N__4962\,
            I => \N__4953\
        );

    \I__1113\ : InMux
    port map (
            O => \N__4959\,
            I => \N__4950\
        );

    \I__1112\ : Sp12to4
    port map (
            O => \N__4956\,
            I => \N__4943\
        );

    \I__1111\ : Sp12to4
    port map (
            O => \N__4953\,
            I => \N__4943\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__4950\,
            I => \N__4943\
        );

    \I__1109\ : Odrv12
    port map (
            O => \N__4943\,
            I => \A_c_6\
        );

    \I__1108\ : CascadeMux
    port map (
            O => \N__4940\,
            I => \N__4930\
        );

    \I__1107\ : InMux
    port map (
            O => \N__4939\,
            I => \N__4925\
        );

    \I__1106\ : CascadeMux
    port map (
            O => \N__4938\,
            I => \N__4920\
        );

    \I__1105\ : CascadeMux
    port map (
            O => \N__4937\,
            I => \N__4917\
        );

    \I__1104\ : InMux
    port map (
            O => \N__4936\,
            I => \N__4914\
        );

    \I__1103\ : InMux
    port map (
            O => \N__4935\,
            I => \N__4911\
        );

    \I__1102\ : InMux
    port map (
            O => \N__4934\,
            I => \N__4908\
        );

    \I__1101\ : InMux
    port map (
            O => \N__4933\,
            I => \N__4903\
        );

    \I__1100\ : InMux
    port map (
            O => \N__4930\,
            I => \N__4900\
        );

    \I__1099\ : InMux
    port map (
            O => \N__4929\,
            I => \N__4897\
        );

    \I__1098\ : InMux
    port map (
            O => \N__4928\,
            I => \N__4894\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__4925\,
            I => \N__4891\
        );

    \I__1096\ : InMux
    port map (
            O => \N__4924\,
            I => \N__4888\
        );

    \I__1095\ : InMux
    port map (
            O => \N__4923\,
            I => \N__4884\
        );

    \I__1094\ : InMux
    port map (
            O => \N__4920\,
            I => \N__4881\
        );

    \I__1093\ : InMux
    port map (
            O => \N__4917\,
            I => \N__4878\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__4914\,
            I => \N__4871\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__4911\,
            I => \N__4871\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__4908\,
            I => \N__4871\
        );

    \I__1089\ : InMux
    port map (
            O => \N__4907\,
            I => \N__4868\
        );

    \I__1088\ : InMux
    port map (
            O => \N__4906\,
            I => \N__4865\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__4903\,
            I => \N__4858\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__4900\,
            I => \N__4858\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__4897\,
            I => \N__4858\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__4894\,
            I => \N__4855\
        );

    \I__1083\ : Span4Mux_h
    port map (
            O => \N__4891\,
            I => \N__4852\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__4888\,
            I => \N__4849\
        );

    \I__1081\ : InMux
    port map (
            O => \N__4887\,
            I => \N__4846\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__4884\,
            I => \N__4839\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__4881\,
            I => \N__4839\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__4878\,
            I => \N__4839\
        );

    \I__1077\ : Span4Mux_v
    port map (
            O => \N__4871\,
            I => \N__4836\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__4868\,
            I => \N__4831\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__4865\,
            I => \N__4831\
        );

    \I__1074\ : Span4Mux_h
    port map (
            O => \N__4858\,
            I => \N__4827\
        );

    \I__1073\ : Span4Mux_h
    port map (
            O => \N__4855\,
            I => \N__4824\
        );

    \I__1072\ : Span4Mux_h
    port map (
            O => \N__4852\,
            I => \N__4817\
        );

    \I__1071\ : Span4Mux_v
    port map (
            O => \N__4849\,
            I => \N__4817\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__4846\,
            I => \N__4817\
        );

    \I__1069\ : Span4Mux_v
    port map (
            O => \N__4839\,
            I => \N__4814\
        );

    \I__1068\ : Span4Mux_h
    port map (
            O => \N__4836\,
            I => \N__4809\
        );

    \I__1067\ : Span4Mux_v
    port map (
            O => \N__4831\,
            I => \N__4809\
        );

    \I__1066\ : InMux
    port map (
            O => \N__4830\,
            I => \N__4806\
        );

    \I__1065\ : Span4Mux_h
    port map (
            O => \N__4827\,
            I => \N__4803\
        );

    \I__1064\ : Span4Mux_h
    port map (
            O => \N__4824\,
            I => \N__4800\
        );

    \I__1063\ : Span4Mux_v
    port map (
            O => \N__4817\,
            I => \N__4797\
        );

    \I__1062\ : Sp12to4
    port map (
            O => \N__4814\,
            I => \N__4790\
        );

    \I__1061\ : Sp12to4
    port map (
            O => \N__4809\,
            I => \N__4790\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__4806\,
            I => \N__4790\
        );

    \I__1059\ : Span4Mux_h
    port map (
            O => \N__4803\,
            I => \N__4785\
        );

    \I__1058\ : Span4Mux_v
    port map (
            O => \N__4800\,
            I => \N__4785\
        );

    \I__1057\ : Span4Mux_h
    port map (
            O => \N__4797\,
            I => \N__4782\
        );

    \I__1056\ : Span12Mux_h
    port map (
            O => \N__4790\,
            I => \N__4779\
        );

    \I__1055\ : Odrv4
    port map (
            O => \N__4785\,
            I => \A_c_1\
        );

    \I__1054\ : Odrv4
    port map (
            O => \N__4782\,
            I => \A_c_1\
        );

    \I__1053\ : Odrv12
    port map (
            O => \N__4779\,
            I => \A_c_1\
        );

    \I__1052\ : IoInMux
    port map (
            O => \N__4772\,
            I => \N__4769\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__4769\,
            I => \N__4766\
        );

    \I__1050\ : Span12Mux_s3_v
    port map (
            O => \N__4766\,
            I => \N__4763\
        );

    \I__1049\ : Odrv12
    port map (
            O => \N__4763\,
            I => \UNGATED_RA_1\
        );

    \I__1048\ : CascadeMux
    port map (
            O => \N__4760\,
            I => \N__4755\
        );

    \I__1047\ : CascadeMux
    port map (
            O => \N__4759\,
            I => \N__4752\
        );

    \I__1046\ : CascadeMux
    port map (
            O => \N__4758\,
            I => \N__4745\
        );

    \I__1045\ : InMux
    port map (
            O => \N__4755\,
            I => \N__4738\
        );

    \I__1044\ : InMux
    port map (
            O => \N__4752\,
            I => \N__4735\
        );

    \I__1043\ : InMux
    port map (
            O => \N__4751\,
            I => \N__4732\
        );

    \I__1042\ : InMux
    port map (
            O => \N__4750\,
            I => \N__4729\
        );

    \I__1041\ : InMux
    port map (
            O => \N__4749\,
            I => \N__4726\
        );

    \I__1040\ : InMux
    port map (
            O => \N__4748\,
            I => \N__4723\
        );

    \I__1039\ : InMux
    port map (
            O => \N__4745\,
            I => \N__4720\
        );

    \I__1038\ : InMux
    port map (
            O => \N__4744\,
            I => \N__4717\
        );

    \I__1037\ : InMux
    port map (
            O => \N__4743\,
            I => \N__4714\
        );

    \I__1036\ : InMux
    port map (
            O => \N__4742\,
            I => \N__4710\
        );

    \I__1035\ : InMux
    port map (
            O => \N__4741\,
            I => \N__4707\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__4738\,
            I => \N__4699\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__4735\,
            I => \N__4699\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__4732\,
            I => \N__4699\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__4729\,
            I => \N__4688\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__4726\,
            I => \N__4688\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__4723\,
            I => \N__4688\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__4720\,
            I => \N__4688\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__4717\,
            I => \N__4688\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__4714\,
            I => \N__4685\
        );

    \I__1025\ : InMux
    port map (
            O => \N__4713\,
            I => \N__4682\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__4710\,
            I => \N__4679\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__4707\,
            I => \N__4676\
        );

    \I__1022\ : InMux
    port map (
            O => \N__4706\,
            I => \N__4673\
        );

    \I__1021\ : Span4Mux_v
    port map (
            O => \N__4699\,
            I => \N__4667\
        );

    \I__1020\ : Span4Mux_v
    port map (
            O => \N__4688\,
            I => \N__4667\
        );

    \I__1019\ : Span4Mux_v
    port map (
            O => \N__4685\,
            I => \N__4662\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__4682\,
            I => \N__4662\
        );

    \I__1017\ : Span4Mux_h
    port map (
            O => \N__4679\,
            I => \N__4655\
        );

    \I__1016\ : Span4Mux_v
    port map (
            O => \N__4676\,
            I => \N__4655\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__4673\,
            I => \N__4655\
        );

    \I__1014\ : InMux
    port map (
            O => \N__4672\,
            I => \N__4651\
        );

    \I__1013\ : Span4Mux_h
    port map (
            O => \N__4667\,
            I => \N__4646\
        );

    \I__1012\ : Span4Mux_v
    port map (
            O => \N__4662\,
            I => \N__4646\
        );

    \I__1011\ : Span4Mux_v
    port map (
            O => \N__4655\,
            I => \N__4643\
        );

    \I__1010\ : InMux
    port map (
            O => \N__4654\,
            I => \N__4640\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__4651\,
            I => \N__4637\
        );

    \I__1008\ : Sp12to4
    port map (
            O => \N__4646\,
            I => \N__4630\
        );

    \I__1007\ : Sp12to4
    port map (
            O => \N__4643\,
            I => \N__4630\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__4640\,
            I => \N__4630\
        );

    \I__1005\ : Span12Mux_h
    port map (
            O => \N__4637\,
            I => \N__4627\
        );

    \I__1004\ : Span12Mux_h
    port map (
            O => \N__4630\,
            I => \N__4624\
        );

    \I__1003\ : Odrv12
    port map (
            O => \N__4627\,
            I => \A_c_2\
        );

    \I__1002\ : Odrv12
    port map (
            O => \N__4624\,
            I => \A_c_2\
        );

    \I__1001\ : InMux
    port map (
            O => \N__4619\,
            I => \N__4613\
        );

    \I__1000\ : InMux
    port map (
            O => \N__4618\,
            I => \N__4610\
        );

    \I__999\ : InMux
    port map (
            O => \N__4617\,
            I => \N__4605\
        );

    \I__998\ : InMux
    port map (
            O => \N__4616\,
            I => \N__4605\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__4613\,
            I => \N__4601\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__4610\,
            I => \N__4596\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__4605\,
            I => \N__4596\
        );

    \I__994\ : InMux
    port map (
            O => \N__4604\,
            I => \N__4593\
        );

    \I__993\ : Span4Mux_h
    port map (
            O => \N__4601\,
            I => \N__4584\
        );

    \I__992\ : Span4Mux_v
    port map (
            O => \N__4596\,
            I => \N__4584\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__4593\,
            I => \N__4584\
        );

    \I__990\ : InMux
    port map (
            O => \N__4592\,
            I => \N__4581\
        );

    \I__989\ : InMux
    port map (
            O => \N__4591\,
            I => \N__4578\
        );

    \I__988\ : Span4Mux_h
    port map (
            O => \N__4584\,
            I => \N__4570\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__4581\,
            I => \N__4570\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__4578\,
            I => \N__4570\
        );

    \I__985\ : InMux
    port map (
            O => \N__4577\,
            I => \N__4567\
        );

    \I__984\ : Odrv4
    port map (
            O => \N__4570\,
            I => \U_MMU_RA.MMU_RA_MUX.D_RAS_N\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__4567\,
            I => \U_MMU_RA.MMU_RA_MUX.D_RAS_N\
        );

    \I__982\ : InMux
    port map (
            O => \N__4562\,
            I => \N__4558\
        );

    \I__981\ : CascadeMux
    port map (
            O => \N__4561\,
            I => \N__4551\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__4558\,
            I => \N__4546\
        );

    \I__979\ : InMux
    port map (
            O => \N__4557\,
            I => \N__4543\
        );

    \I__978\ : InMux
    port map (
            O => \N__4556\,
            I => \N__4538\
        );

    \I__977\ : InMux
    port map (
            O => \N__4555\,
            I => \N__4538\
        );

    \I__976\ : InMux
    port map (
            O => \N__4554\,
            I => \N__4535\
        );

    \I__975\ : InMux
    port map (
            O => \N__4551\,
            I => \N__4532\
        );

    \I__974\ : InMux
    port map (
            O => \N__4550\,
            I => \N__4529\
        );

    \I__973\ : CascadeMux
    port map (
            O => \N__4549\,
            I => \N__4525\
        );

    \I__972\ : Span4Mux_h
    port map (
            O => \N__4546\,
            I => \N__4522\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__4543\,
            I => \N__4517\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__4538\,
            I => \N__4517\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__4535\,
            I => \N__4512\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__4532\,
            I => \N__4512\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__4529\,
            I => \N__4509\
        );

    \I__966\ : InMux
    port map (
            O => \N__4528\,
            I => \N__4506\
        );

    \I__965\ : InMux
    port map (
            O => \N__4525\,
            I => \N__4503\
        );

    \I__964\ : Span4Mux_h
    port map (
            O => \N__4522\,
            I => \N__4496\
        );

    \I__963\ : Span4Mux_h
    port map (
            O => \N__4517\,
            I => \N__4496\
        );

    \I__962\ : Span4Mux_v
    port map (
            O => \N__4512\,
            I => \N__4491\
        );

    \I__961\ : Span4Mux_h
    port map (
            O => \N__4509\,
            I => \N__4491\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4506\,
            I => \N__4486\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__4503\,
            I => \N__4486\
        );

    \I__958\ : InMux
    port map (
            O => \N__4502\,
            I => \N__4483\
        );

    \I__957\ : InMux
    port map (
            O => \N__4501\,
            I => \N__4480\
        );

    \I__956\ : Span4Mux_v
    port map (
            O => \N__4496\,
            I => \N__4477\
        );

    \I__955\ : Span4Mux_h
    port map (
            O => \N__4491\,
            I => \N__4472\
        );

    \I__954\ : Span4Mux_v
    port map (
            O => \N__4486\,
            I => \N__4472\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__4483\,
            I => \N__4467\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__4480\,
            I => \N__4467\
        );

    \I__951\ : Sp12to4
    port map (
            O => \N__4477\,
            I => \N__4460\
        );

    \I__950\ : Sp12to4
    port map (
            O => \N__4472\,
            I => \N__4460\
        );

    \I__949\ : Span12Mux_h
    port map (
            O => \N__4467\,
            I => \N__4460\
        );

    \I__948\ : Odrv12
    port map (
            O => \N__4460\,
            I => \PRAS_N_c\
        );

    \I__947\ : InMux
    port map (
            O => \N__4457\,
            I => \N__4454\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__4454\,
            I => \N__4450\
        );

    \I__945\ : InMux
    port map (
            O => \N__4453\,
            I => \N__4444\
        );

    \I__944\ : Span4Mux_h
    port map (
            O => \N__4450\,
            I => \N__4441\
        );

    \I__943\ : InMux
    port map (
            O => \N__4449\,
            I => \N__4438\
        );

    \I__942\ : InMux
    port map (
            O => \N__4448\,
            I => \N__4434\
        );

    \I__941\ : InMux
    port map (
            O => \N__4447\,
            I => \N__4431\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__4444\,
            I => \N__4427\
        );

    \I__939\ : Span4Mux_v
    port map (
            O => \N__4441\,
            I => \N__4422\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__4438\,
            I => \N__4422\
        );

    \I__937\ : InMux
    port map (
            O => \N__4437\,
            I => \N__4419\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__4434\,
            I => \N__4416\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__4431\,
            I => \N__4413\
        );

    \I__934\ : InMux
    port map (
            O => \N__4430\,
            I => \N__4410\
        );

    \I__933\ : Span4Mux_h
    port map (
            O => \N__4427\,
            I => \N__4407\
        );

    \I__932\ : Span4Mux_h
    port map (
            O => \N__4422\,
            I => \N__4404\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__4419\,
            I => \N__4401\
        );

    \I__930\ : Span4Mux_h
    port map (
            O => \N__4416\,
            I => \N__4396\
        );

    \I__929\ : Span4Mux_h
    port map (
            O => \N__4413\,
            I => \N__4396\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__4410\,
            I => \N__4393\
        );

    \I__927\ : Span4Mux_v
    port map (
            O => \N__4407\,
            I => \N__4390\
        );

    \I__926\ : Span4Mux_v
    port map (
            O => \N__4404\,
            I => \N__4387\
        );

    \I__925\ : Span4Mux_h
    port map (
            O => \N__4401\,
            I => \N__4384\
        );

    \I__924\ : Span4Mux_v
    port map (
            O => \N__4396\,
            I => \N__4379\
        );

    \I__923\ : Span4Mux_h
    port map (
            O => \N__4393\,
            I => \N__4379\
        );

    \I__922\ : Odrv4
    port map (
            O => \N__4390\,
            I => \A_c_10\
        );

    \I__921\ : Odrv4
    port map (
            O => \N__4387\,
            I => \A_c_10\
        );

    \I__920\ : Odrv4
    port map (
            O => \N__4384\,
            I => \A_c_10\
        );

    \I__919\ : Odrv4
    port map (
            O => \N__4379\,
            I => \A_c_10\
        );

    \I__918\ : IoInMux
    port map (
            O => \N__4370\,
            I => \N__4367\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__4367\,
            I => \N__4364\
        );

    \I__916\ : Span12Mux_s11_v
    port map (
            O => \N__4364\,
            I => \N__4361\
        );

    \I__915\ : Odrv12
    port map (
            O => \N__4361\,
            I => \UNGATED_RA_2\
        );

    \I__914\ : IoInMux
    port map (
            O => \N__4358\,
            I => \N__4355\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__4355\,
            I => \ORA_pad_0AndNet\
        );

    \I__912\ : SRMux
    port map (
            O => \N__4352\,
            I => \N__4349\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__4349\,
            I => \N__4346\
        );

    \I__910\ : Span4Mux_v
    port map (
            O => \N__4346\,
            I => \N__4343\
        );

    \I__909\ : Odrv4
    port map (
            O => \N__4343\,
            I => \U_MMU_RA.MMU_RA_MUX.RA_ENABLE_N_N_215\
        );

    \I__908\ : InMux
    port map (
            O => \N__4340\,
            I => \N__4336\
        );

    \I__907\ : InMux
    port map (
            O => \N__4339\,
            I => \N__4333\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__4336\,
            I => \RA_ENABLE_N\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__4333\,
            I => \RA_ENABLE_N\
        );

    \I__904\ : IoInMux
    port map (
            O => \N__4328\,
            I => \N__4325\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__4325\,
            I => \ORA_pad_3AndNet\
        );

    \I__902\ : IoInMux
    port map (
            O => \N__4322\,
            I => \N__4319\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__4319\,
            I => \ORA_pad_4AndNet\
        );

    \I__900\ : IoInMux
    port map (
            O => \N__4316\,
            I => \N__4313\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__4313\,
            I => \ORA_pad_5AndNet\
        );

    \I__898\ : InMux
    port map (
            O => \N__4310\,
            I => \N__4307\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__4307\,
            I => \ORA_pad_3LegalizeSB_DFFNet\
        );

    \I__896\ : InMux
    port map (
            O => \N__4304\,
            I => \N__4301\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__4301\,
            I => \ORA_pad_4LegalizeSB_DFFNet\
        );

    \I__894\ : InMux
    port map (
            O => \N__4298\,
            I => \N__4295\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__4295\,
            I => \ORA_pad_5LegalizeSB_DFFNet\
        );

    \I__892\ : InMux
    port map (
            O => \N__4292\,
            I => \N__4288\
        );

    \I__891\ : InMux
    port map (
            O => \N__4291\,
            I => \N__4285\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__4288\,
            I => \N__4281\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__4285\,
            I => \N__4278\
        );

    \I__888\ : InMux
    port map (
            O => \N__4284\,
            I => \N__4275\
        );

    \I__887\ : Span4Mux_h
    port map (
            O => \N__4281\,
            I => \N__4272\
        );

    \I__886\ : Span4Mux_h
    port map (
            O => \N__4278\,
            I => \N__4267\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__4275\,
            I => \N__4267\
        );

    \I__884\ : Span4Mux_v
    port map (
            O => \N__4272\,
            I => \N__4261\
        );

    \I__883\ : Span4Mux_h
    port map (
            O => \N__4267\,
            I => \N__4261\
        );

    \I__882\ : InMux
    port map (
            O => \N__4266\,
            I => \N__4258\
        );

    \I__881\ : Sp12to4
    port map (
            O => \N__4261\,
            I => \N__4255\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__4258\,
            I => \N__4252\
        );

    \I__879\ : Odrv12
    port map (
            O => \N__4255\,
            I => \Q3_c\
        );

    \I__878\ : Odrv4
    port map (
            O => \N__4252\,
            I => \Q3_c\
        );

    \I__877\ : CascadeMux
    port map (
            O => \N__4247\,
            I => \N__4241\
        );

    \I__876\ : CascadeMux
    port map (
            O => \N__4246\,
            I => \N__4233\
        );

    \I__875\ : CascadeMux
    port map (
            O => \N__4245\,
            I => \N__4229\
        );

    \I__874\ : CascadeMux
    port map (
            O => \N__4244\,
            I => \N__4226\
        );

    \I__873\ : InMux
    port map (
            O => \N__4241\,
            I => \N__4222\
        );

    \I__872\ : InMux
    port map (
            O => \N__4240\,
            I => \N__4219\
        );

    \I__871\ : InMux
    port map (
            O => \N__4239\,
            I => \N__4216\
        );

    \I__870\ : InMux
    port map (
            O => \N__4238\,
            I => \N__4213\
        );

    \I__869\ : InMux
    port map (
            O => \N__4237\,
            I => \N__4210\
        );

    \I__868\ : InMux
    port map (
            O => \N__4236\,
            I => \N__4207\
        );

    \I__867\ : InMux
    port map (
            O => \N__4233\,
            I => \N__4204\
        );

    \I__866\ : InMux
    port map (
            O => \N__4232\,
            I => \N__4201\
        );

    \I__865\ : InMux
    port map (
            O => \N__4229\,
            I => \N__4198\
        );

    \I__864\ : InMux
    port map (
            O => \N__4226\,
            I => \N__4195\
        );

    \I__863\ : InMux
    port map (
            O => \N__4225\,
            I => \N__4192\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__4222\,
            I => \N__4189\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__4219\,
            I => \N__4186\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__4216\,
            I => \N__4183\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__4213\,
            I => \N__4180\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__4210\,
            I => \N__4177\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__4207\,
            I => \N__4174\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__4204\,
            I => \N__4171\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__4201\,
            I => \N__4167\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__4198\,
            I => \N__4164\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__4195\,
            I => \N__4161\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__4192\,
            I => \N__4158\
        );

    \I__851\ : Glb2LocalMux
    port map (
            O => \N__4189\,
            I => \N__4133\
        );

    \I__850\ : Glb2LocalMux
    port map (
            O => \N__4186\,
            I => \N__4133\
        );

    \I__849\ : Glb2LocalMux
    port map (
            O => \N__4183\,
            I => \N__4133\
        );

    \I__848\ : Glb2LocalMux
    port map (
            O => \N__4180\,
            I => \N__4133\
        );

    \I__847\ : Glb2LocalMux
    port map (
            O => \N__4177\,
            I => \N__4133\
        );

    \I__846\ : Glb2LocalMux
    port map (
            O => \N__4174\,
            I => \N__4133\
        );

    \I__845\ : Glb2LocalMux
    port map (
            O => \N__4171\,
            I => \N__4133\
        );

    \I__844\ : ClkMux
    port map (
            O => \N__4170\,
            I => \N__4133\
        );

    \I__843\ : Glb2LocalMux
    port map (
            O => \N__4167\,
            I => \N__4133\
        );

    \I__842\ : Glb2LocalMux
    port map (
            O => \N__4164\,
            I => \N__4133\
        );

    \I__841\ : Glb2LocalMux
    port map (
            O => \N__4161\,
            I => \N__4133\
        );

    \I__840\ : Glb2LocalMux
    port map (
            O => \N__4158\,
            I => \N__4133\
        );

    \I__839\ : GlobalMux
    port map (
            O => \N__4133\,
            I => \N__4130\
        );

    \I__838\ : gio2CtrlBuf
    port map (
            O => \N__4130\,
            I => \PHI_0_c\
        );

    \I__837\ : InMux
    port map (
            O => \N__4127\,
            I => \N__4124\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__4124\,
            I => \U_ADDR_DECODER.n9\
        );

    \I__835\ : InMux
    port map (
            O => \N__4121\,
            I => \N__4118\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__4118\,
            I => \U_MMU_MPON.n13\
        );

    \I__833\ : CascadeMux
    port map (
            O => \N__4115\,
            I => \N__4111\
        );

    \I__832\ : CascadeMux
    port map (
            O => \N__4114\,
            I => \N__4107\
        );

    \I__831\ : InMux
    port map (
            O => \N__4111\,
            I => \N__4104\
        );

    \I__830\ : InMux
    port map (
            O => \N__4110\,
            I => \N__4101\
        );

    \I__829\ : InMux
    port map (
            O => \N__4107\,
            I => \N__4098\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__4104\,
            I => \N__4095\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__4101\,
            I => \N__4091\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__4098\,
            I => \N__4088\
        );

    \I__825\ : Span4Mux_h
    port map (
            O => \N__4095\,
            I => \N__4085\
        );

    \I__824\ : CascadeMux
    port map (
            O => \N__4094\,
            I => \N__4081\
        );

    \I__823\ : Span4Mux_h
    port map (
            O => \N__4091\,
            I => \N__4078\
        );

    \I__822\ : Span4Mux_h
    port map (
            O => \N__4088\,
            I => \N__4075\
        );

    \I__821\ : Span4Mux_v
    port map (
            O => \N__4085\,
            I => \N__4072\
        );

    \I__820\ : InMux
    port map (
            O => \N__4084\,
            I => \N__4069\
        );

    \I__819\ : InMux
    port map (
            O => \N__4081\,
            I => \N__4066\
        );

    \I__818\ : Span4Mux_v
    port map (
            O => \N__4078\,
            I => \N__4063\
        );

    \I__817\ : Span4Mux_v
    port map (
            O => \N__4075\,
            I => \N__4060\
        );

    \I__816\ : Sp12to4
    port map (
            O => \N__4072\,
            I => \N__4053\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__4069\,
            I => \N__4053\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__4066\,
            I => \N__4053\
        );

    \I__813\ : Odrv4
    port map (
            O => \N__4063\,
            I => \A_c_8\
        );

    \I__812\ : Odrv4
    port map (
            O => \N__4060\,
            I => \A_c_8\
        );

    \I__811\ : Odrv12
    port map (
            O => \N__4053\,
            I => \A_c_8\
        );

    \I__810\ : InMux
    port map (
            O => \N__4046\,
            I => \N__4043\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__4043\,
            I => \N__4039\
        );

    \I__808\ : InMux
    port map (
            O => \N__4042\,
            I => \N__4036\
        );

    \I__807\ : Span4Mux_v
    port map (
            O => \N__4039\,
            I => \N__4033\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__4036\,
            I => \N__4030\
        );

    \I__805\ : Odrv4
    port map (
            O => \N__4033\,
            I => n626
        );

    \I__804\ : Odrv4
    port map (
            O => \N__4030\,
            I => n626
        );

    \I__803\ : InMux
    port map (
            O => \N__4025\,
            I => \N__4019\
        );

    \I__802\ : InMux
    port map (
            O => \N__4024\,
            I => \N__4019\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__4019\,
            I => \U_MMU_MPON.M5_2\
        );

    \I__800\ : InMux
    port map (
            O => \N__4016\,
            I => \N__4012\
        );

    \I__799\ : InMux
    port map (
            O => \N__4015\,
            I => \N__4009\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__4012\,
            I => \U_MMU_MPON.M5_7\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__4009\,
            I => \U_MMU_MPON.M5_7\
        );

    \I__796\ : InMux
    port map (
            O => \N__4004\,
            I => \N__4001\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__4001\,
            I => \U_MMU_MPON.DELTA_01XX_N\
        );

    \I__794\ : InMux
    port map (
            O => \N__3998\,
            I => \N__3995\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__3995\,
            I => n2523
        );

    \I__792\ : InMux
    port map (
            O => \N__3992\,
            I => \N__3988\
        );

    \I__791\ : InMux
    port map (
            O => \N__3991\,
            I => \N__3985\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__3988\,
            I => \N__3981\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__3985\,
            I => \N__3975\
        );

    \I__788\ : InMux
    port map (
            O => \N__3984\,
            I => \N__3971\
        );

    \I__787\ : Span4Mux_v
    port map (
            O => \N__3981\,
            I => \N__3968\
        );

    \I__786\ : InMux
    port map (
            O => \N__3980\,
            I => \N__3965\
        );

    \I__785\ : InMux
    port map (
            O => \N__3979\,
            I => \N__3960\
        );

    \I__784\ : InMux
    port map (
            O => \N__3978\,
            I => \N__3960\
        );

    \I__783\ : Span4Mux_h
    port map (
            O => \N__3975\,
            I => \N__3957\
        );

    \I__782\ : InMux
    port map (
            O => \N__3974\,
            I => \N__3954\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__3971\,
            I => \N__3951\
        );

    \I__780\ : Span4Mux_h
    port map (
            O => \N__3968\,
            I => \N__3942\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__3965\,
            I => \N__3942\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__3960\,
            I => \N__3942\
        );

    \I__777\ : Span4Mux_h
    port map (
            O => \N__3957\,
            I => \N__3936\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__3954\,
            I => \N__3936\
        );

    \I__775\ : Span4Mux_v
    port map (
            O => \N__3951\,
            I => \N__3933\
        );

    \I__774\ : InMux
    port map (
            O => \N__3950\,
            I => \N__3930\
        );

    \I__773\ : InMux
    port map (
            O => \N__3949\,
            I => \N__3927\
        );

    \I__772\ : Span4Mux_v
    port map (
            O => \N__3942\,
            I => \N__3924\
        );

    \I__771\ : InMux
    port map (
            O => \N__3941\,
            I => \N__3921\
        );

    \I__770\ : Span4Mux_v
    port map (
            O => \N__3936\,
            I => \N__3918\
        );

    \I__769\ : Sp12to4
    port map (
            O => \N__3933\,
            I => \N__3907\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__3930\,
            I => \N__3907\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__3927\,
            I => \N__3907\
        );

    \I__766\ : Sp12to4
    port map (
            O => \N__3924\,
            I => \N__3907\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__3921\,
            I => \N__3907\
        );

    \I__764\ : Sp12to4
    port map (
            O => \N__3918\,
            I => \N__3902\
        );

    \I__763\ : Span12Mux_h
    port map (
            O => \N__3907\,
            I => \N__3902\
        );

    \I__762\ : Odrv12
    port map (
            O => \N__3902\,
            I => \R_W_N_c\
        );

    \I__761\ : CascadeMux
    port map (
            O => \N__3899\,
            I => \n2523_cascade_\
        );

    \I__760\ : InMux
    port map (
            O => \N__3896\,
            I => \N__3893\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__3893\,
            I => \U_ADDR_DECODER.n7\
        );

    \I__758\ : InMux
    port map (
            O => \N__3890\,
            I => \N__3887\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__3887\,
            I => n906
        );

    \I__756\ : CascadeMux
    port map (
            O => \N__3884\,
            I => \n953_cascade_\
        );

    \I__755\ : ClkMux
    port map (
            O => \N__3881\,
            I => \N__3877\
        );

    \I__754\ : ClkMux
    port map (
            O => \N__3880\,
            I => \N__3874\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__3877\,
            I => \N__3871\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__3874\,
            I => \N__3867\
        );

    \I__751\ : Span4Mux_v
    port map (
            O => \N__3871\,
            I => \N__3864\
        );

    \I__750\ : ClkMux
    port map (
            O => \N__3870\,
            I => \N__3861\
        );

    \I__749\ : Span4Mux_v
    port map (
            O => \N__3867\,
            I => \N__3858\
        );

    \I__748\ : Span4Mux_h
    port map (
            O => \N__3864\,
            I => \N__3855\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__3861\,
            I => \N__3852\
        );

    \I__746\ : Odrv4
    port map (
            O => \N__3858\,
            I => \DEV0_N\
        );

    \I__745\ : Odrv4
    port map (
            O => \N__3855\,
            I => \DEV0_N\
        );

    \I__744\ : Odrv12
    port map (
            O => \N__3852\,
            I => \DEV0_N\
        );

    \I__743\ : InMux
    port map (
            O => \N__3845\,
            I => \N__3842\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__3842\,
            I => n953
        );

    \I__741\ : CascadeMux
    port map (
            O => \N__3839\,
            I => \ENABLE_N_cascade_\
        );

    \I__740\ : InMux
    port map (
            O => \N__3836\,
            I => \N__3833\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__3833\,
            I => \N__3830\
        );

    \I__738\ : Odrv4
    port map (
            O => \N__3830\,
            I => n912
        );

    \I__737\ : CascadeMux
    port map (
            O => \N__3827\,
            I => \N__3822\
        );

    \I__736\ : InMux
    port map (
            O => \N__3826\,
            I => \N__3818\
        );

    \I__735\ : InMux
    port map (
            O => \N__3825\,
            I => \N__3815\
        );

    \I__734\ : InMux
    port map (
            O => \N__3822\,
            I => \N__3812\
        );

    \I__733\ : InMux
    port map (
            O => \N__3821\,
            I => \N__3809\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__3818\,
            I => \MC0XX_N\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__3815\,
            I => \MC0XX_N\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__3812\,
            I => \MC0XX_N\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__3809\,
            I => \MC0XX_N\
        );

    \I__728\ : CascadeMux
    port map (
            O => \N__3800\,
            I => \N__3796\
        );

    \I__727\ : CascadeMux
    port map (
            O => \N__3799\,
            I => \N__3792\
        );

    \I__726\ : InMux
    port map (
            O => \N__3796\,
            I => \N__3789\
        );

    \I__725\ : CascadeMux
    port map (
            O => \N__3795\,
            I => \N__3784\
        );

    \I__724\ : InMux
    port map (
            O => \N__3792\,
            I => \N__3780\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__3789\,
            I => \N__3777\
        );

    \I__722\ : InMux
    port map (
            O => \N__3788\,
            I => \N__3774\
        );

    \I__721\ : InMux
    port map (
            O => \N__3787\,
            I => \N__3771\
        );

    \I__720\ : InMux
    port map (
            O => \N__3784\,
            I => \N__3768\
        );

    \I__719\ : CascadeMux
    port map (
            O => \N__3783\,
            I => \N__3765\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__3780\,
            I => \N__3762\
        );

    \I__717\ : Span4Mux_v
    port map (
            O => \N__3777\,
            I => \N__3754\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__3774\,
            I => \N__3754\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__3771\,
            I => \N__3754\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__3768\,
            I => \N__3751\
        );

    \I__713\ : InMux
    port map (
            O => \N__3765\,
            I => \N__3748\
        );

    \I__712\ : Span4Mux_h
    port map (
            O => \N__3762\,
            I => \N__3745\
        );

    \I__711\ : InMux
    port map (
            O => \N__3761\,
            I => \N__3742\
        );

    \I__710\ : Span4Mux_h
    port map (
            O => \N__3754\,
            I => \N__3739\
        );

    \I__709\ : Span4Mux_h
    port map (
            O => \N__3751\,
            I => \N__3736\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__3748\,
            I => \N__3733\
        );

    \I__707\ : Span4Mux_v
    port map (
            O => \N__3745\,
            I => \N__3730\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__3742\,
            I => \N__3727\
        );

    \I__705\ : Span4Mux_v
    port map (
            O => \N__3739\,
            I => \N__3724\
        );

    \I__704\ : Span4Mux_v
    port map (
            O => \N__3736\,
            I => \N__3719\
        );

    \I__703\ : Span4Mux_h
    port map (
            O => \N__3733\,
            I => \N__3719\
        );

    \I__702\ : Sp12to4
    port map (
            O => \N__3730\,
            I => \N__3714\
        );

    \I__701\ : Span12Mux_h
    port map (
            O => \N__3727\,
            I => \N__3714\
        );

    \I__700\ : Odrv4
    port map (
            O => \N__3724\,
            I => \A_c_7\
        );

    \I__699\ : Odrv4
    port map (
            O => \N__3719\,
            I => \A_c_7\
        );

    \I__698\ : Odrv12
    port map (
            O => \N__3714\,
            I => \A_c_7\
        );

    \I__697\ : InMux
    port map (
            O => \N__3707\,
            I => \N__3704\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__3704\,
            I => \N__3700\
        );

    \I__695\ : InMux
    port map (
            O => \N__3703\,
            I => \N__3697\
        );

    \I__694\ : Span4Mux_v
    port map (
            O => \N__3700\,
            I => \N__3693\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__3697\,
            I => \N__3690\
        );

    \I__692\ : CascadeMux
    port map (
            O => \N__3696\,
            I => \N__3687\
        );

    \I__691\ : Span4Mux_h
    port map (
            O => \N__3693\,
            I => \N__3682\
        );

    \I__690\ : Span4Mux_v
    port map (
            O => \N__3690\,
            I => \N__3682\
        );

    \I__689\ : InMux
    port map (
            O => \N__3687\,
            I => \N__3679\
        );

    \I__688\ : Odrv4
    port map (
            O => \N__3682\,
            I => \U_ADDR_DECODER.n44\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__3679\,
            I => \U_ADDR_DECODER.n44\
        );

    \I__686\ : InMux
    port map (
            O => \N__3674\,
            I => \N__3671\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__3671\,
            I => \N__3668\
        );

    \I__684\ : Span12Mux_s10_h
    port map (
            O => \N__3668\,
            I => \N__3665\
        );

    \I__683\ : Span12Mux_v
    port map (
            O => \N__3665\,
            I => \N__3662\
        );

    \I__682\ : Odrv12
    port map (
            O => \N__3662\,
            I => \MD7_ENABLE_N_N_6\
        );

    \I__681\ : CascadeMux
    port map (
            O => \N__3659\,
            I => \N__3655\
        );

    \I__680\ : InMux
    port map (
            O => \N__3658\,
            I => \N__3651\
        );

    \I__679\ : InMux
    port map (
            O => \N__3655\,
            I => \N__3644\
        );

    \I__678\ : InMux
    port map (
            O => \N__3654\,
            I => \N__3644\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__3651\,
            I => \N__3641\
        );

    \I__676\ : InMux
    port map (
            O => \N__3650\,
            I => \N__3636\
        );

    \I__675\ : InMux
    port map (
            O => \N__3649\,
            I => \N__3636\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__3644\,
            I => \N__3632\
        );

    \I__673\ : Span4Mux_v
    port map (
            O => \N__3641\,
            I => \N__3627\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__3636\,
            I => \N__3627\
        );

    \I__671\ : InMux
    port map (
            O => \N__3635\,
            I => \N__3624\
        );

    \I__670\ : Span4Mux_h
    port map (
            O => \N__3632\,
            I => \N__3621\
        );

    \I__669\ : Span4Mux_h
    port map (
            O => \N__3627\,
            I => \N__3616\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__3624\,
            I => \N__3616\
        );

    \I__667\ : Span4Mux_v
    port map (
            O => \N__3621\,
            I => \N__3613\
        );

    \I__666\ : Span4Mux_h
    port map (
            O => \N__3616\,
            I => \N__3610\
        );

    \I__665\ : Odrv4
    port map (
            O => \N__3613\,
            I => \A_c_13\
        );

    \I__664\ : Odrv4
    port map (
            O => \N__3610\,
            I => \A_c_13\
        );

    \I__663\ : InMux
    port map (
            O => \N__3605\,
            I => \N__3599\
        );

    \I__662\ : InMux
    port map (
            O => \N__3604\,
            I => \N__3596\
        );

    \I__661\ : InMux
    port map (
            O => \N__3603\,
            I => \N__3593\
        );

    \I__660\ : InMux
    port map (
            O => \N__3602\,
            I => \N__3589\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__3599\,
            I => \N__3582\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__3596\,
            I => \N__3582\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__3593\,
            I => \N__3582\
        );

    \I__656\ : InMux
    port map (
            O => \N__3592\,
            I => \N__3579\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__3589\,
            I => \N__3576\
        );

    \I__654\ : Span4Mux_v
    port map (
            O => \N__3582\,
            I => \N__3570\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__3579\,
            I => \N__3570\
        );

    \I__652\ : Span4Mux_v
    port map (
            O => \N__3576\,
            I => \N__3567\
        );

    \I__651\ : InMux
    port map (
            O => \N__3575\,
            I => \N__3564\
        );

    \I__650\ : Span4Mux_v
    port map (
            O => \N__3570\,
            I => \N__3561\
        );

    \I__649\ : Sp12to4
    port map (
            O => \N__3567\,
            I => \N__3556\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__3564\,
            I => \N__3556\
        );

    \I__647\ : Span4Mux_h
    port map (
            O => \N__3561\,
            I => \N__3553\
        );

    \I__646\ : Span12Mux_h
    port map (
            O => \N__3556\,
            I => \N__3550\
        );

    \I__645\ : Odrv4
    port map (
            O => \N__3553\,
            I => \A_c_5\
        );

    \I__644\ : Odrv12
    port map (
            O => \N__3550\,
            I => \A_c_5\
        );

    \I__643\ : IoInMux
    port map (
            O => \N__3545\,
            I => \N__3542\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__3542\,
            I => \N__3539\
        );

    \I__641\ : Span4Mux_s1_v
    port map (
            O => \N__3539\,
            I => \N__3536\
        );

    \I__640\ : Span4Mux_v
    port map (
            O => \N__3536\,
            I => \N__3533\
        );

    \I__639\ : Span4Mux_v
    port map (
            O => \N__3533\,
            I => \N__3530\
        );

    \I__638\ : Odrv4
    port map (
            O => \N__3530\,
            I => \UNGATED_RA_5\
        );

    \I__637\ : InMux
    port map (
            O => \N__3527\,
            I => \N__3521\
        );

    \I__636\ : InMux
    port map (
            O => \N__3526\,
            I => \N__3518\
        );

    \I__635\ : InMux
    port map (
            O => \N__3525\,
            I => \N__3514\
        );

    \I__634\ : InMux
    port map (
            O => \N__3524\,
            I => \N__3511\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__3521\,
            I => \N__3505\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__3518\,
            I => \N__3505\
        );

    \I__631\ : InMux
    port map (
            O => \N__3517\,
            I => \N__3502\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__3514\,
            I => \N__3497\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__3511\,
            I => \N__3497\
        );

    \I__628\ : InMux
    port map (
            O => \N__3510\,
            I => \N__3494\
        );

    \I__627\ : Span4Mux_v
    port map (
            O => \N__3505\,
            I => \N__3491\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__3502\,
            I => \N__3484\
        );

    \I__625\ : Span4Mux_v
    port map (
            O => \N__3497\,
            I => \N__3484\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__3494\,
            I => \N__3484\
        );

    \I__623\ : Sp12to4
    port map (
            O => \N__3491\,
            I => \N__3479\
        );

    \I__622\ : Sp12to4
    port map (
            O => \N__3484\,
            I => \N__3479\
        );

    \I__621\ : Span12Mux_h
    port map (
            O => \N__3479\,
            I => \N__3476\
        );

    \I__620\ : Odrv12
    port map (
            O => \N__3476\,
            I => \A_c_4\
        );

    \I__619\ : CascadeMux
    port map (
            O => \N__3473\,
            I => \MC0XX_N_cascade_\
        );

    \I__618\ : InMux
    port map (
            O => \N__3470\,
            I => \N__3467\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__3467\,
            I => n2576
        );

    \I__616\ : CascadeMux
    port map (
            O => \N__3464\,
            I => \n1226_cascade_\
        );

    \I__615\ : InMux
    port map (
            O => \N__3461\,
            I => \N__3455\
        );

    \I__614\ : InMux
    port map (
            O => \N__3460\,
            I => \N__3455\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__3455\,
            I => \N__3452\
        );

    \I__612\ : Span4Mux_v
    port map (
            O => \N__3452\,
            I => \N__3449\
        );

    \I__611\ : Odrv4
    port map (
            O => \N__3449\,
            I => \LATCHED_MC05X_N\
        );

    \I__610\ : InMux
    port map (
            O => \N__3446\,
            I => \N__3443\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__3443\,
            I => n933
        );

    \I__608\ : InMux
    port map (
            O => \N__3440\,
            I => \N__3437\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__3437\,
            I => \UMMU_INTERNALS.n2580\
        );

    \I__606\ : InMux
    port map (
            O => \N__3434\,
            I => \N__3431\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__3431\,
            I => n2520
        );

    \I__604\ : InMux
    port map (
            O => \N__3428\,
            I => \N__3425\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__3425\,
            I => \N__3422\
        );

    \I__602\ : Span4Mux_v
    port map (
            O => \N__3422\,
            I => \N__3419\
        );

    \I__601\ : Odrv4
    port map (
            O => \N__3419\,
            I => \MA12_N_209\
        );

    \I__600\ : CascadeMux
    port map (
            O => \N__3416\,
            I => \U_MMU_RA.MMU_RA_MUX.COMBINED_RAS_N_cascade_\
        );

    \I__599\ : InMux
    port map (
            O => \N__3413\,
            I => \N__3406\
        );

    \I__598\ : InMux
    port map (
            O => \N__3412\,
            I => \N__3403\
        );

    \I__597\ : InMux
    port map (
            O => \N__3411\,
            I => \N__3398\
        );

    \I__596\ : InMux
    port map (
            O => \N__3410\,
            I => \N__3398\
        );

    \I__595\ : InMux
    port map (
            O => \N__3409\,
            I => \N__3395\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__3406\,
            I => \N__3392\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__3403\,
            I => \N__3388\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__3398\,
            I => \N__3385\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__3395\,
            I => \N__3382\
        );

    \I__590\ : Span4Mux_h
    port map (
            O => \N__3392\,
            I => \N__3379\
        );

    \I__589\ : InMux
    port map (
            O => \N__3391\,
            I => \N__3372\
        );

    \I__588\ : Span4Mux_v
    port map (
            O => \N__3388\,
            I => \N__3367\
        );

    \I__587\ : Span4Mux_h
    port map (
            O => \N__3385\,
            I => \N__3367\
        );

    \I__586\ : Span4Mux_h
    port map (
            O => \N__3382\,
            I => \N__3364\
        );

    \I__585\ : Span4Mux_h
    port map (
            O => \N__3379\,
            I => \N__3361\
        );

    \I__584\ : InMux
    port map (
            O => \N__3378\,
            I => \N__3354\
        );

    \I__583\ : InMux
    port map (
            O => \N__3377\,
            I => \N__3354\
        );

    \I__582\ : InMux
    port map (
            O => \N__3376\,
            I => \N__3354\
        );

    \I__581\ : InMux
    port map (
            O => \N__3375\,
            I => \N__3351\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__3372\,
            I => \N__3348\
        );

    \I__579\ : Span4Mux_h
    port map (
            O => \N__3367\,
            I => \N__3345\
        );

    \I__578\ : Span4Mux_v
    port map (
            O => \N__3364\,
            I => \N__3342\
        );

    \I__577\ : Sp12to4
    port map (
            O => \N__3361\,
            I => \N__3335\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__3354\,
            I => \N__3335\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__3351\,
            I => \N__3335\
        );

    \I__574\ : Span4Mux_h
    port map (
            O => \N__3348\,
            I => \N__3332\
        );

    \I__573\ : Odrv4
    port map (
            O => \N__3345\,
            I => \A_c_12\
        );

    \I__572\ : Odrv4
    port map (
            O => \N__3342\,
            I => \A_c_12\
        );

    \I__571\ : Odrv12
    port map (
            O => \N__3335\,
            I => \A_c_12\
        );

    \I__570\ : Odrv4
    port map (
            O => \N__3332\,
            I => \A_c_12\
        );

    \I__569\ : IoInMux
    port map (
            O => \N__3323\,
            I => \N__3320\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__3320\,
            I => \N__3317\
        );

    \I__567\ : Span4Mux_s3_v
    port map (
            O => \N__3317\,
            I => \N__3314\
        );

    \I__566\ : Span4Mux_v
    port map (
            O => \N__3314\,
            I => \N__3311\
        );

    \I__565\ : Span4Mux_v
    port map (
            O => \N__3311\,
            I => \N__3308\
        );

    \I__564\ : Odrv4
    port map (
            O => \N__3308\,
            I => \UNGATED_RA_4\
        );

    \I__563\ : InMux
    port map (
            O => \N__3305\,
            I => \N__3302\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__3302\,
            I => \U_MMU_RA.MMU_RA_MUX.U_DRAM_HOLD_TIME.PRAS_N_SHIFT_REGISTER_2\
        );

    \I__561\ : ClkMux
    port map (
            O => \N__3299\,
            I => \N__3275\
        );

    \I__560\ : ClkMux
    port map (
            O => \N__3298\,
            I => \N__3275\
        );

    \I__559\ : ClkMux
    port map (
            O => \N__3297\,
            I => \N__3275\
        );

    \I__558\ : ClkMux
    port map (
            O => \N__3296\,
            I => \N__3275\
        );

    \I__557\ : ClkMux
    port map (
            O => \N__3295\,
            I => \N__3275\
        );

    \I__556\ : ClkMux
    port map (
            O => \N__3294\,
            I => \N__3275\
        );

    \I__555\ : ClkMux
    port map (
            O => \N__3293\,
            I => \N__3275\
        );

    \I__554\ : ClkMux
    port map (
            O => \N__3292\,
            I => \N__3275\
        );

    \I__553\ : GlobalMux
    port map (
            O => \N__3275\,
            I => \DELAY_CLK\
        );

    \I__552\ : InMux
    port map (
            O => \N__3272\,
            I => \N__3269\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__3269\,
            I => \U_ADDR_DECODER.S_0XXX_N\
        );

    \I__550\ : IoInMux
    port map (
            O => \N__3266\,
            I => \N__3263\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3263\,
            I => \N__3260\
        );

    \I__548\ : Span4Mux_s1_v
    port map (
            O => \N__3260\,
            I => \N__3257\
        );

    \I__547\ : Span4Mux_v
    port map (
            O => \N__3257\,
            I => \N__3254\
        );

    \I__546\ : Span4Mux_v
    port map (
            O => \N__3254\,
            I => \N__3251\
        );

    \I__545\ : Odrv4
    port map (
            O => \N__3251\,
            I => \UNGATED_RA_7\
        );

    \I__544\ : InMux
    port map (
            O => \N__3248\,
            I => \N__3245\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__3245\,
            I => \U_MMU_RA.MMU_RA_MUX.U_DRAM_HOLD_TIME.PRAS_N_SHIFT_REGISTER_0\
        );

    \I__542\ : InMux
    port map (
            O => \N__3242\,
            I => \N__3239\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__3239\,
            I => \U_MMU_RA.MMU_RA_MUX.U_DRAM_HOLD_TIME.PRAS_N_SHIFT_REGISTER_1\
        );

    \I__540\ : InMux
    port map (
            O => \N__3236\,
            I => \N__3232\
        );

    \I__539\ : CascadeMux
    port map (
            O => \N__3235\,
            I => \N__3226\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__3232\,
            I => \N__3223\
        );

    \I__537\ : InMux
    port map (
            O => \N__3231\,
            I => \N__3218\
        );

    \I__536\ : InMux
    port map (
            O => \N__3230\,
            I => \N__3218\
        );

    \I__535\ : InMux
    port map (
            O => \N__3229\,
            I => \N__3215\
        );

    \I__534\ : InMux
    port map (
            O => \N__3226\,
            I => \N__3212\
        );

    \I__533\ : Span4Mux_h
    port map (
            O => \N__3223\,
            I => \N__3208\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__3218\,
            I => \N__3205\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__3215\,
            I => \N__3200\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__3212\,
            I => \N__3200\
        );

    \I__529\ : InMux
    port map (
            O => \N__3211\,
            I => \N__3197\
        );

    \I__528\ : Span4Mux_h
    port map (
            O => \N__3208\,
            I => \N__3194\
        );

    \I__527\ : Span4Mux_h
    port map (
            O => \N__3205\,
            I => \N__3191\
        );

    \I__526\ : Span4Mux_h
    port map (
            O => \N__3200\,
            I => \N__3186\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__3197\,
            I => \N__3186\
        );

    \I__524\ : Sp12to4
    port map (
            O => \N__3194\,
            I => \N__3183\
        );

    \I__523\ : Span4Mux_v
    port map (
            O => \N__3191\,
            I => \N__3180\
        );

    \I__522\ : Span4Mux_h
    port map (
            O => \N__3186\,
            I => \N__3177\
        );

    \I__521\ : Odrv12
    port map (
            O => \N__3183\,
            I => \A_c_14\
        );

    \I__520\ : Odrv4
    port map (
            O => \N__3180\,
            I => \A_c_14\
        );

    \I__519\ : Odrv4
    port map (
            O => \N__3177\,
            I => \A_c_14\
        );

    \I__518\ : InMux
    port map (
            O => \N__3170\,
            I => \N__3167\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__3167\,
            I => \N__3164\
        );

    \I__516\ : Span4Mux_v
    port map (
            O => \N__3164\,
            I => \N__3157\
        );

    \I__515\ : InMux
    port map (
            O => \N__3163\,
            I => \N__3152\
        );

    \I__514\ : InMux
    port map (
            O => \N__3162\,
            I => \N__3152\
        );

    \I__513\ : InMux
    port map (
            O => \N__3161\,
            I => \N__3147\
        );

    \I__512\ : InMux
    port map (
            O => \N__3160\,
            I => \N__3147\
        );

    \I__511\ : Span4Mux_v
    port map (
            O => \N__3157\,
            I => \N__3141\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__3152\,
            I => \N__3141\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__3147\,
            I => \N__3138\
        );

    \I__508\ : InMux
    port map (
            O => \N__3146\,
            I => \N__3135\
        );

    \I__507\ : Span4Mux_v
    port map (
            O => \N__3141\,
            I => \N__3132\
        );

    \I__506\ : Span4Mux_v
    port map (
            O => \N__3138\,
            I => \N__3127\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__3135\,
            I => \N__3127\
        );

    \I__504\ : Span4Mux_h
    port map (
            O => \N__3132\,
            I => \N__3122\
        );

    \I__503\ : Span4Mux_v
    port map (
            O => \N__3127\,
            I => \N__3122\
        );

    \I__502\ : Span4Mux_h
    port map (
            O => \N__3122\,
            I => \N__3119\
        );

    \I__501\ : Odrv4
    port map (
            O => \N__3119\,
            I => \A_c_15\
        );

    \I__500\ : InMux
    port map (
            O => \N__3116\,
            I => \N__3113\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__3113\,
            I => \U_MMU_MPON.n2521\
        );

    \I__498\ : CascadeMux
    port map (
            O => \N__3110\,
            I => \U_MMU_MPON.n2602_cascade_\
        );

    \I__497\ : InMux
    port map (
            O => \N__3107\,
            I => \N__3103\
        );

    \I__496\ : InMux
    port map (
            O => \N__3106\,
            I => \N__3100\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__3103\,
            I => \N__3097\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__3100\,
            I => \N__3094\
        );

    \I__493\ : Odrv12
    port map (
            O => \N__3097\,
            I => \U_ADDR_DECODER.MC0XX_N_N_20\
        );

    \I__492\ : Odrv4
    port map (
            O => \N__3094\,
            I => \U_ADDR_DECODER.MC0XX_N_N_20\
        );

    \I__491\ : InMux
    port map (
            O => \N__3089\,
            I => \N__3083\
        );

    \I__490\ : InMux
    port map (
            O => \N__3088\,
            I => \N__3083\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__3083\,
            I => \PENIO_N\
        );

    \I__488\ : CascadeMux
    port map (
            O => \N__3080\,
            I => \PENIO_N_cascade_\
        );

    \I__487\ : InMux
    port map (
            O => \N__3077\,
            I => \N__3074\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__3074\,
            I => \N__3071\
        );

    \I__485\ : Odrv4
    port map (
            O => \N__3071\,
            I => \U_MMU_MD7.n4\
        );

    \I__484\ : CascadeMux
    port map (
            O => \N__3068\,
            I => \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.n2570_cascade_\
        );

    \I__483\ : CascadeMux
    port map (
            O => \N__3065\,
            I => \N__3062\
        );

    \I__482\ : InMux
    port map (
            O => \N__3062\,
            I => \N__3059\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__3059\,
            I => \N__3055\
        );

    \I__480\ : InMux
    port map (
            O => \N__3058\,
            I => \N__3052\
        );

    \I__479\ : Span4Mux_h
    port map (
            O => \N__3055\,
            I => \N__3048\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__3052\,
            I => \N__3045\
        );

    \I__477\ : InMux
    port map (
            O => \N__3051\,
            I => \N__3042\
        );

    \I__476\ : Odrv4
    port map (
            O => \N__3048\,
            I => \EN80VID\
        );

    \I__475\ : Odrv4
    port map (
            O => \N__3045\,
            I => \EN80VID\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__3042\,
            I => \EN80VID\
        );

    \I__473\ : InMux
    port map (
            O => \N__3035\,
            I => \N__3032\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__3032\,
            I => \N__3029\
        );

    \I__471\ : Odrv4
    port map (
            O => \N__3029\,
            I => n927
        );

    \I__470\ : InMux
    port map (
            O => \N__3026\,
            I => \N__3023\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__3023\,
            I => \N__3019\
        );

    \I__468\ : InMux
    port map (
            O => \N__3022\,
            I => \N__3016\
        );

    \I__467\ : Odrv12
    port map (
            O => \N__3019\,
            I => \C8_FXX\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__3016\,
            I => \C8_FXX\
        );

    \I__465\ : CascadeMux
    port map (
            O => \N__3011\,
            I => \n927_cascade_\
        );

    \I__464\ : CascadeMux
    port map (
            O => \N__3008\,
            I => \UMMU_INTERNALS.n2616_cascade_\
        );

    \I__463\ : InMux
    port map (
            O => \N__3005\,
            I => \N__3002\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__3002\,
            I => \N__2999\
        );

    \I__461\ : Odrv4
    port map (
            O => \N__2999\,
            I => \UMMU_INTERNALS.n2622\
        );

    \I__460\ : IoInMux
    port map (
            O => \N__2996\,
            I => \N__2993\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__2993\,
            I => \N__2990\
        );

    \I__458\ : Span12Mux_s1_v
    port map (
            O => \N__2990\,
            I => \N__2987\
        );

    \I__457\ : Odrv12
    port map (
            O => \N__2987\,
            I => \UNGATED_RA_6\
        );

    \I__456\ : IoInMux
    port map (
            O => \N__2984\,
            I => \N__2981\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__2981\,
            I => \N__2978\
        );

    \I__454\ : Span12Mux_s5_v
    port map (
            O => \N__2978\,
            I => \N__2975\
        );

    \I__453\ : Odrv12
    port map (
            O => \N__2975\,
            I => \KBD_N_c\
        );

    \I__452\ : InMux
    port map (
            O => \N__2972\,
            I => \N__2969\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__2969\,
            I => \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.n938\
        );

    \I__450\ : InMux
    port map (
            O => \N__2966\,
            I => \N__2963\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__2963\,
            I => \N__2957\
        );

    \I__448\ : InMux
    port map (
            O => \N__2962\,
            I => \N__2950\
        );

    \I__447\ : InMux
    port map (
            O => \N__2961\,
            I => \N__2950\
        );

    \I__446\ : InMux
    port map (
            O => \N__2960\,
            I => \N__2950\
        );

    \I__445\ : Span4Mux_v
    port map (
            O => \N__2957\,
            I => \N__2945\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__2950\,
            I => \N__2942\
        );

    \I__443\ : InMux
    port map (
            O => \N__2949\,
            I => \N__2939\
        );

    \I__442\ : InMux
    port map (
            O => \N__2948\,
            I => \N__2936\
        );

    \I__441\ : Odrv4
    port map (
            O => \N__2945\,
            I => \DXXX_N_N_13\
        );

    \I__440\ : Odrv4
    port map (
            O => \N__2942\,
            I => \DXXX_N_N_13\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__2939\,
            I => \DXXX_N_N_13\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__2936\,
            I => \DXXX_N_N_13\
        );

    \I__437\ : InMux
    port map (
            O => \N__2927\,
            I => \N__2924\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__2924\,
            I => \BANK1\
        );

    \I__435\ : IoInMux
    port map (
            O => \N__2921\,
            I => \N__2918\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__2918\,
            I => \ORA_pad_6AndNet\
        );

    \I__433\ : IoInMux
    port map (
            O => \N__2915\,
            I => \N__2912\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__2912\,
            I => \ORA_pad_7AndNet\
        );

    \I__431\ : IoInMux
    port map (
            O => \N__2909\,
            I => \N__2906\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__2906\,
            I => \KBD_N_padLegalizeSB_DFFNet\
        );

    \I__429\ : InMux
    port map (
            O => \N__2903\,
            I => \N__2900\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__2900\,
            I => \ORA_pad_6LegalizeSB_DFFNet\
        );

    \I__427\ : InMux
    port map (
            O => \N__2897\,
            I => \N__2894\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__2894\,
            I => \ORA_pad_7LegalizeSB_DFFNet\
        );

    \I__425\ : InMux
    port map (
            O => \N__2891\,
            I => \N__2885\
        );

    \I__424\ : InMux
    port map (
            O => \N__2890\,
            I => \N__2885\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__2885\,
            I => \N__2882\
        );

    \I__422\ : Span4Mux_v
    port map (
            O => \N__2882\,
            I => \N__2879\
        );

    \I__421\ : Odrv4
    port map (
            O => \N__2879\,
            I => \CENROM1\
        );

    \I__420\ : InMux
    port map (
            O => \N__2876\,
            I => \N__2873\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__2873\,
            I => \U_MMU_RA.MMU_RA_MUX.U_DRAM_HOLD_TIME.Q3_SHIFT_REGISTER_0\
        );

    \I__418\ : InMux
    port map (
            O => \N__2870\,
            I => \N__2867\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__2867\,
            I => \U_MMU_RA.MMU_RA_MUX.U_DRAM_HOLD_TIME.Q3_SHIFT_REGISTER_1\
        );

    \I__416\ : InMux
    port map (
            O => \N__2864\,
            I => \N__2861\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__2861\,
            I => \N__2858\
        );

    \I__414\ : Odrv4
    port map (
            O => \N__2858\,
            I => n2584
        );

    \I__413\ : InMux
    port map (
            O => \N__2855\,
            I => \N__2852\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__2852\,
            I => \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.n937\
        );

    \I__411\ : CascadeMux
    port map (
            O => \N__2849\,
            I => \N__2846\
        );

    \I__410\ : InMux
    port map (
            O => \N__2846\,
            I => \N__2843\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__2843\,
            I => \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.n2532\
        );

    \I__408\ : CascadeMux
    port map (
            O => \N__2840\,
            I => \ALTSTKZP_cascade_\
        );

    \I__407\ : InMux
    port map (
            O => \N__2837\,
            I => \N__2834\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__2834\,
            I => \N__2830\
        );

    \I__405\ : InMux
    port map (
            O => \N__2833\,
            I => \N__2827\
        );

    \I__404\ : Odrv4
    port map (
            O => \N__2830\,
            I => \INTC300_N\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__2827\,
            I => \INTC300_N\
        );

    \I__402\ : InMux
    port map (
            O => \N__2822\,
            I => \N__2819\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__2819\,
            I => \U_MMU_MD7.n5\
        );

    \I__400\ : InMux
    port map (
            O => \N__2816\,
            I => \N__2813\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__2813\,
            I => \N__2808\
        );

    \I__398\ : InMux
    port map (
            O => \N__2812\,
            I => \N__2805\
        );

    \I__397\ : InMux
    port map (
            O => \N__2811\,
            I => \N__2802\
        );

    \I__396\ : Odrv4
    port map (
            O => \N__2808\,
            I => \FLG1\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__2805\,
            I => \FLG1\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__2802\,
            I => \FLG1\
        );

    \I__393\ : InMux
    port map (
            O => \N__2795\,
            I => \N__2791\
        );

    \I__392\ : InMux
    port map (
            O => \N__2794\,
            I => \N__2788\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__2791\,
            I => \ALTSTKZP\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__2788\,
            I => \ALTSTKZP\
        );

    \I__389\ : CascadeMux
    port map (
            O => \N__2783\,
            I => \SELMB_N_N_137_cascade_\
        );

    \I__388\ : InMux
    port map (
            O => \N__2780\,
            I => \N__2777\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__2777\,
            I => \N__2774\
        );

    \I__386\ : Span4Mux_h
    port map (
            O => \N__2774\,
            I => \N__2771\
        );

    \I__385\ : Odrv4
    port map (
            O => \N__2771\,
            I => \D_FXXX\
        );

    \I__384\ : InMux
    port map (
            O => \N__2768\,
            I => \N__2765\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__2765\,
            I => \N__2762\
        );

    \I__382\ : Odrv4
    port map (
            O => \N__2762\,
            I => \U_MMU_SELMB.SELMB_N_N_136\
        );

    \I__381\ : InMux
    port map (
            O => \N__2759\,
            I => \N__2756\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__2756\,
            I => \U_MMU_MD7.n2710\
        );

    \I__379\ : IoInMux
    port map (
            O => \N__2753\,
            I => \N__2750\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__2750\,
            I => \N__2747\
        );

    \I__377\ : IoSpan4Mux
    port map (
            O => \N__2747\,
            I => \N__2744\
        );

    \I__376\ : Span4Mux_s2_v
    port map (
            O => \N__2744\,
            I => \N__2741\
        );

    \I__375\ : Sp12to4
    port map (
            O => \N__2741\,
            I => \N__2738\
        );

    \I__374\ : Span12Mux_v
    port map (
            O => \N__2738\,
            I => \N__2735\
        );

    \I__373\ : Odrv12
    port map (
            O => \N__2735\,
            I => \UNGATED_MD7\
        );

    \I__372\ : InMux
    port map (
            O => \N__2732\,
            I => \N__2729\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__2729\,
            I => \U_MMU_MD7.n2707\
        );

    \I__370\ : InMux
    port map (
            O => \N__2726\,
            I => \N__2723\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__2723\,
            I => \BANK2\
        );

    \I__368\ : InMux
    port map (
            O => \N__2720\,
            I => \N__2717\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__2717\,
            I => \N__2714\
        );

    \I__366\ : Odrv12
    port map (
            O => \N__2714\,
            I => \RDROM\
        );

    \I__365\ : CascadeMux
    port map (
            O => \N__2711\,
            I => \INTC300_N_cascade_\
        );

    \I__364\ : InMux
    port map (
            O => \N__2708\,
            I => \N__2702\
        );

    \I__363\ : InMux
    port map (
            O => \N__2707\,
            I => \N__2702\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__2702\,
            I => \N__2698\
        );

    \I__361\ : InMux
    port map (
            O => \N__2701\,
            I => \N__2695\
        );

    \I__360\ : Odrv12
    port map (
            O => \N__2698\,
            I => \INTC3ACC_N_N_175\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__2695\,
            I => \INTC3ACC_N_N_175\
        );

    \I__358\ : ClkMux
    port map (
            O => \N__2690\,
            I => \N__2687\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__2687\,
            I => \N__2684\
        );

    \I__356\ : Span4Mux_v
    port map (
            O => \N__2684\,
            I => \N__2681\
        );

    \I__355\ : Span4Mux_h
    port map (
            O => \N__2681\,
            I => \N__2678\
        );

    \I__354\ : Odrv4
    port map (
            O => \N__2678\,
            I => \U_MMU_RA.MMU_RA_MUX.D_Q3\
        );

    \I__353\ : CascadeMux
    port map (
            O => \N__2675\,
            I => \UMMU_INTERNALS.n1605_cascade_\
        );

    \I__352\ : InMux
    port map (
            O => \N__2672\,
            I => \N__2665\
        );

    \I__351\ : InMux
    port map (
            O => \N__2671\,
            I => \N__2665\
        );

    \I__350\ : InMux
    port map (
            O => \N__2670\,
            I => \N__2662\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__2665\,
            I => \INTC8EN\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__2662\,
            I => \INTC8EN\
        );

    \I__347\ : CascadeMux
    port map (
            O => \N__2657\,
            I => \N__2654\
        );

    \I__346\ : InMux
    port map (
            O => \N__2654\,
            I => \N__2651\
        );

    \I__345\ : LocalMux
    port map (
            O => \N__2651\,
            I => \U_MMU_HOLD_TIME.SHIFT_REGISTER_1\
        );

    \I__344\ : InMux
    port map (
            O => \N__2648\,
            I => \N__2645\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__2645\,
            I => \U_MMU_HOLD_TIME.SHIFT_REGISTER_0\
        );

    \I__342\ : InMux
    port map (
            O => \N__2642\,
            I => \N__2639\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__2639\,
            I => \N__2636\
        );

    \I__340\ : Odrv4
    port map (
            O => \N__2636\,
            I => n2596
        );

    \I__339\ : InMux
    port map (
            O => \N__2633\,
            I => \N__2630\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__2630\,
            I => n911
        );

    \I__337\ : InMux
    port map (
            O => \N__2627\,
            I => \N__2624\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2624\,
            I => \RDRAM\
        );

    \I__335\ : CascadeMux
    port map (
            O => \N__2621\,
            I => \U_MMU_MD7.n2658_cascade_\
        );

    \I__334\ : InMux
    port map (
            O => \N__2618\,
            I => \N__2615\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__2615\,
            I => \U_MMU_MD7.n2\
        );

    \I__332\ : InMux
    port map (
            O => \N__2612\,
            I => \N__2609\
        );

    \I__331\ : LocalMux
    port map (
            O => \N__2609\,
            I => \U_MMU_SELMB.n2572\
        );

    \I__330\ : InMux
    port map (
            O => \N__2606\,
            I => \N__2603\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__2603\,
            I => \U_MMU_SELMB.n2610\
        );

    \I__328\ : CascadeMux
    port map (
            O => \N__2600\,
            I => \HIRES_cascade_\
        );

    \I__327\ : InMux
    port map (
            O => \N__2597\,
            I => \N__2594\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__2594\,
            I => \N__2591\
        );

    \I__325\ : Odrv4
    port map (
            O => \N__2591\,
            I => \WRPROT\
        );

    \I__324\ : CascadeMux
    port map (
            O => \N__2588\,
            I => \N__2585\
        );

    \I__323\ : InMux
    port map (
            O => \N__2585\,
            I => \N__2581\
        );

    \I__322\ : InMux
    port map (
            O => \N__2584\,
            I => \N__2578\
        );

    \I__321\ : LocalMux
    port map (
            O => \N__2581\,
            I => \U_MMU_SOFT_SWITCHES_C08X.OUT_FST_ACC\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__2578\,
            I => \U_MMU_SOFT_SWITCHES_C08X.OUT_FST_ACC\
        );

    \I__319\ : CascadeMux
    port map (
            O => \N__2573\,
            I => \N__2569\
        );

    \I__318\ : InMux
    port map (
            O => \N__2572\,
            I => \N__2564\
        );

    \I__317\ : InMux
    port map (
            O => \N__2569\,
            I => \N__2564\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__2564\,
            I => \U_MMU_SOFT_SWITCHES_C08X.OUT_WREN\
        );

    \I__315\ : InMux
    port map (
            O => \N__2561\,
            I => \N__2558\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__2558\,
            I => \N__2555\
        );

    \I__313\ : Odrv4
    port map (
            O => \N__2555\,
            I => \U_MMU_SELMB.n2516\
        );

    \I__312\ : CascadeMux
    port map (
            O => \N__2552\,
            I => \N__2549\
        );

    \I__311\ : InMux
    port map (
            O => \N__2549\,
            I => \N__2545\
        );

    \I__310\ : InMux
    port map (
            O => \N__2548\,
            I => \N__2542\
        );

    \I__309\ : LocalMux
    port map (
            O => \N__2545\,
            I => \PG2\
        );

    \I__308\ : LocalMux
    port map (
            O => \N__2542\,
            I => \PG2\
        );

    \I__307\ : InMux
    port map (
            O => \N__2537\,
            I => \N__2533\
        );

    \I__306\ : InMux
    port map (
            O => \N__2536\,
            I => \N__2530\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__2533\,
            I => \N__2525\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__2530\,
            I => \N__2525\
        );

    \I__303\ : Span4Mux_v
    port map (
            O => \N__2525\,
            I => \N__2522\
        );

    \I__302\ : Odrv4
    port map (
            O => \N__2522\,
            I => \SELMB_N\
        );

    \I__301\ : CascadeMux
    port map (
            O => \N__2519\,
            I => \N__2515\
        );

    \I__300\ : InMux
    port map (
            O => \N__2518\,
            I => \N__2512\
        );

    \I__299\ : InMux
    port map (
            O => \N__2515\,
            I => \N__2508\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__2512\,
            I => \N__2505\
        );

    \I__297\ : InMux
    port map (
            O => \N__2511\,
            I => \N__2502\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__2508\,
            I => \N__2499\
        );

    \I__295\ : Odrv4
    port map (
            O => \N__2505\,
            I => \D_PHI_0\
        );

    \I__294\ : LocalMux
    port map (
            O => \N__2502\,
            I => \D_PHI_0\
        );

    \I__293\ : Odrv12
    port map (
            O => \N__2499\,
            I => \D_PHI_0\
        );

    \I__292\ : InMux
    port map (
            O => \N__2492\,
            I => \N__2489\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__2489\,
            I => \INTC8ACC\
        );

    \I__290\ : CascadeMux
    port map (
            O => \N__2486\,
            I => \CXXX_cascade_\
        );

    \I__289\ : InMux
    port map (
            O => \N__2483\,
            I => \N__2480\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__2480\,
            I => n966
        );

    \I__287\ : InMux
    port map (
            O => \N__2477\,
            I => \N__2474\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__2474\,
            I => \CXXX\
        );

    \I__285\ : InMux
    port map (
            O => \N__2471\,
            I => \N__2468\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__2468\,
            I => \U_MMU_ROMEN.n7\
        );

    \I__283\ : CascadeMux
    port map (
            O => \N__2465\,
            I => \N__2462\
        );

    \I__282\ : InMux
    port map (
            O => \N__2462\,
            I => \N__2459\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__2459\,
            I => \U_MMU_ROMEN.n4\
        );

    \I__280\ : IoInMux
    port map (
            O => \N__2456\,
            I => \N__2453\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__2453\,
            I => \N__2450\
        );

    \I__278\ : Span4Mux_s3_v
    port map (
            O => \N__2450\,
            I => \N__2447\
        );

    \I__277\ : Sp12to4
    port map (
            O => \N__2447\,
            I => \N__2444\
        );

    \I__276\ : Span12Mux_s9_h
    port map (
            O => \N__2444\,
            I => \N__2441\
        );

    \I__275\ : Odrv12
    port map (
            O => \N__2441\,
            I => \ROMEN1_N_INT\
        );

    \I__274\ : InMux
    port map (
            O => \N__2438\,
            I => \N__2430\
        );

    \I__273\ : InMux
    port map (
            O => \N__2437\,
            I => \N__2430\
        );

    \I__272\ : InMux
    port map (
            O => \N__2436\,
            I => \N__2427\
        );

    \I__271\ : InMux
    port map (
            O => \N__2435\,
            I => \N__2424\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__2430\,
            I => \N__2421\
        );

    \I__269\ : LocalMux
    port map (
            O => \N__2427\,
            I => \N__2418\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__2424\,
            I => \N__2415\
        );

    \I__267\ : Span4Mux_h
    port map (
            O => \N__2421\,
            I => \N__2412\
        );

    \I__266\ : Span4Mux_h
    port map (
            O => \N__2418\,
            I => \N__2407\
        );

    \I__265\ : Span4Mux_h
    port map (
            O => \N__2415\,
            I => \N__2407\
        );

    \I__264\ : Sp12to4
    port map (
            O => \N__2412\,
            I => \N__2404\
        );

    \I__263\ : Span4Mux_v
    port map (
            O => \N__2407\,
            I => \N__2401\
        );

    \I__262\ : Odrv12
    port map (
            O => \N__2404\,
            I => \INH_N_c\
        );

    \I__261\ : Odrv4
    port map (
            O => \N__2401\,
            I => \INH_N_c\
        );

    \I__260\ : IoInMux
    port map (
            O => \N__2396\,
            I => \N__2393\
        );

    \I__259\ : LocalMux
    port map (
            O => \N__2393\,
            I => \N__2390\
        );

    \I__258\ : Span12Mux_s7_v
    port map (
            O => \N__2390\,
            I => \N__2386\
        );

    \I__257\ : InMux
    port map (
            O => \N__2389\,
            I => \N__2383\
        );

    \I__256\ : Odrv12
    port map (
            O => \N__2386\,
            I => \CXXXOUT_c\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__2383\,
            I => \CXXXOUT_c\
        );

    \I__254\ : InMux
    port map (
            O => \N__2378\,
            I => \N__2375\
        );

    \I__253\ : LocalMux
    port map (
            O => \N__2375\,
            I => \N__2372\
        );

    \I__252\ : Odrv12
    port map (
            O => \N__2372\,
            I => \U_ADDR_DECODER.n2654\
        );

    \I__251\ : IoInMux
    port map (
            O => \N__2369\,
            I => \N__2366\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__2366\,
            I => \N__2363\
        );

    \I__249\ : Span12Mux_s0_v
    port map (
            O => \N__2363\,
            I => \N__2360\
        );

    \I__248\ : Odrv12
    port map (
            O => \N__2360\,
            I => \EN80_N_c\
        );

    \I__247\ : InMux
    port map (
            O => \N__2357\,
            I => \N__2353\
        );

    \I__246\ : InMux
    port map (
            O => \N__2356\,
            I => \N__2350\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__2353\,
            I => \N__2345\
        );

    \I__244\ : LocalMux
    port map (
            O => \N__2350\,
            I => \N__2345\
        );

    \I__243\ : Odrv4
    port map (
            O => \N__2345\,
            I => n907
        );

    \I__242\ : IoInMux
    port map (
            O => \N__2342\,
            I => \N__2339\
        );

    \I__241\ : LocalMux
    port map (
            O => \N__2339\,
            I => \N__2336\
        );

    \I__240\ : IoSpan4Mux
    port map (
            O => \N__2336\,
            I => \N__2333\
        );

    \I__239\ : Sp12to4
    port map (
            O => \N__2333\,
            I => \N__2330\
        );

    \I__238\ : Odrv12
    port map (
            O => \N__2330\,
            I => \CASEN_N_c\
        );

    \I__237\ : InMux
    port map (
            O => \N__2327\,
            I => \N__2324\
        );

    \I__236\ : LocalMux
    port map (
            O => \N__2324\,
            I => \HIRES\
        );

    \I__235\ : InMux
    port map (
            O => \N__2321\,
            I => \N__2318\
        );

    \I__234\ : LocalMux
    port map (
            O => \N__2318\,
            I => \N__2314\
        );

    \I__233\ : InMux
    port map (
            O => \N__2317\,
            I => \N__2311\
        );

    \I__232\ : Odrv4
    port map (
            O => \N__2314\,
            I => \FXXX_N_N_8\
        );

    \I__231\ : LocalMux
    port map (
            O => \N__2311\,
            I => \FXXX_N_N_8\
        );

    \I__230\ : CascadeMux
    port map (
            O => \N__2306\,
            I => \D_FXXX_cascade_\
        );

    \I__229\ : CascadeMux
    port map (
            O => \N__2303\,
            I => \N__2300\
        );

    \I__228\ : InMux
    port map (
            O => \N__2300\,
            I => \N__2295\
        );

    \I__227\ : InMux
    port map (
            O => \N__2299\,
            I => \N__2292\
        );

    \I__226\ : InMux
    port map (
            O => \N__2298\,
            I => \N__2289\
        );

    \I__225\ : LocalMux
    port map (
            O => \N__2295\,
            I => \D2_6_N_148\
        );

    \I__224\ : LocalMux
    port map (
            O => \N__2292\,
            I => \D2_6_N_148\
        );

    \I__223\ : LocalMux
    port map (
            O => \N__2289\,
            I => \D2_6_N_148\
        );

    \I__222\ : CascadeMux
    port map (
            O => \N__2282\,
            I => \C8_FXX_cascade_\
        );

    \I__221\ : InMux
    port map (
            O => \N__2279\,
            I => \N__2276\
        );

    \I__220\ : LocalMux
    port map (
            O => \N__2276\,
            I => \N__2273\
        );

    \I__219\ : Odrv12
    port map (
            O => \N__2273\,
            I => \DMA_N_c\
        );

    \I__218\ : IoInMux
    port map (
            O => \N__2270\,
            I => \N__2267\
        );

    \I__217\ : LocalMux
    port map (
            O => \N__2267\,
            I => \N__2264\
        );

    \I__216\ : Span4Mux_s3_v
    port map (
            O => \N__2264\,
            I => \N__2261\
        );

    \I__215\ : Span4Mux_v
    port map (
            O => \N__2261\,
            I => \N__2258\
        );

    \I__214\ : Span4Mux_v
    port map (
            O => \N__2258\,
            I => \N__2255\
        );

    \I__213\ : Odrv4
    port map (
            O => \N__2255\,
            I => \R_W_N_245_INT\
        );

    \I__212\ : IoInMux
    port map (
            O => \N__2252\,
            I => \N__2249\
        );

    \I__211\ : LocalMux
    port map (
            O => \N__2249\,
            I => \U_MD7AndNet\
        );

    \I__210\ : InMux
    port map (
            O => \N__2246\,
            I => \N__2243\
        );

    \I__209\ : LocalMux
    port map (
            O => \N__2243\,
            I => \U_MD7LegalizeSB_DFFNet\
        );

    \I__208\ : IoInMux
    port map (
            O => \N__2240\,
            I => \N__2237\
        );

    \I__207\ : LocalMux
    port map (
            O => \N__2237\,
            I => \U_ROMEN1_NLegalizeSB_DFFNet\
        );

    \I__206\ : IoInMux
    port map (
            O => \N__2234\,
            I => \N__2231\
        );

    \I__205\ : LocalMux
    port map (
            O => \N__2231\,
            I => \N__2228\
        );

    \I__204\ : Span12Mux_s4_v
    port map (
            O => \N__2228\,
            I => \N__2225\
        );

    \I__203\ : Odrv12
    port map (
            O => \N__2225\,
            I => \ROMEN2_N_c\
        );

    \I__202\ : IoInMux
    port map (
            O => \N__2222\,
            I => \N__2219\
        );

    \I__201\ : LocalMux
    port map (
            O => \N__2219\,
            I => \CASEN_N_padLegalizeSB_DFFNet\
        );

    \I__200\ : IoInMux
    port map (
            O => \N__2216\,
            I => \N__2213\
        );

    \I__199\ : LocalMux
    port map (
            O => \N__2213\,
            I => \CXXXOUT_padLegalizeSB_DFFNet\
        );

    \I__198\ : IoInMux
    port map (
            O => \N__2210\,
            I => \N__2207\
        );

    \I__197\ : LocalMux
    port map (
            O => \N__2207\,
            I => \EN80_N_padLegalizeSB_DFFNet\
        );

    \I__196\ : IoInMux
    port map (
            O => \N__2204\,
            I => \N__2201\
        );

    \I__195\ : LocalMux
    port map (
            O => \N__2201\,
            I => \ROMEN2_N_padLegalizeSB_DFFNet\
        );

    \I__194\ : InMux
    port map (
            O => \N__2198\,
            I => \N__2194\
        );

    \I__193\ : InMux
    port map (
            O => \N__2197\,
            I => \N__2191\
        );

    \I__192\ : LocalMux
    port map (
            O => \N__2194\,
            I => \CONSTANT_ONE_NET\
        );

    \I__191\ : LocalMux
    port map (
            O => \N__2191\,
            I => \CONSTANT_ONE_NET\
        );

    \I__190\ : IoInMux
    port map (
            O => \N__2186\,
            I => \N__2183\
        );

    \I__189\ : LocalMux
    port map (
            O => \N__2183\,
            I => \U_R_W_N_245LegalizeSB_DFFNet\
        );

    \INVU_MMU_RA.MMU_RA_MUX.RA_ENABLE_N_22C\ : INV
    port map (
            O => \INVU_MMU_RA.MMU_RA_MUX.RA_ENABLE_N_22C_net\,
            I => \N__2690\
        );

    \INVU_MMU_SOFT_SWITCHES_C08X.RDROM_31C\ : INV
    port map (
            O => \INVU_MMU_SOFT_SWITCHES_C08X.RDROM_31C_net\,
            I => \N__3880\
        );

    \INVU_MMU_SOFT_SWITCHES_C08X.BANK2_30C\ : INV
    port map (
            O => \INVU_MMU_SOFT_SWITCHES_C08X.BANK2_30C_net\,
            I => \N__3881\
        );

    \INVU_MMU_SOFT_SWITCHES_C08X.OUT_FST_ACC_27C\ : INV
    port map (
            O => \INVU_MMU_SOFT_SWITCHES_C08X.OUT_FST_ACC_27C_net\,
            I => \N__3870\
        );

    \internalOscilator\ : SMCCLK
    port map (
            CLK => \internalOscilatorOutputNet\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \U_DELAY_OSCILLATOR.U_SB_HFOSC\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b00"
        )
    port map (
            CLKHFPU => \N__2198\,
            CLKHFEN => \N__2197\,
            CLKHF => \DELAY_CLK\
        );

    \U_ROMEN1_N\ : SB_IO_OD
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PACKAGEPIN => ROMEN1_N,
            INPUTCLK => '0',
            OUTPUTENABLE => \N__2240\,
            LATCHINPUTVALUE => '0',
            DOUT1 => \GNDG0\,
            DIN1 => OPEN,
            OUTPUTCLK => '0',
            DOUT0 => \N__2456\,
            DIN0 => OPEN,
            CLOCKENABLE => '0'
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \U_MD7\ : SB_IO_OD
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PACKAGEPIN => MD7,
            INPUTCLK => '0',
            OUTPUTENABLE => \N__2252\,
            LATCHINPUTVALUE => '0',
            DOUT1 => \GNDG0\,
            DIN1 => OPEN,
            OUTPUTCLK => '0',
            DOUT0 => \N__2753\,
            DIN0 => OPEN,
            CLOCKENABLE => '0'
        );

    \U_R_W_N_245\ : SB_IO_OD
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PACKAGEPIN => R_W_N_245,
            INPUTCLK => '0',
            OUTPUTENABLE => \N__2186\,
            LATCHINPUTVALUE => '0',
            DOUT1 => \GNDG0\,
            DIN1 => OPEN,
            OUTPUTCLK => '0',
            DOUT0 => \N__2270\,
            DIN0 => OPEN,
            CLOCKENABLE => '0'
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_1_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_R_W_N_245LegalizeSB_DFF_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U_R_W_N_245LegalizeSB_DFFNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5762\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_ADDR_DECODER.i1_4_lut_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001110000"
        )
    port map (
            in0 => \N__2378\,
            in1 => \N__3974\,
            in2 => \N__4247\,
            in3 => \N__2279\,
            lcout => \R_W_N_245_INT\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MD7AndLUT4_LC_5_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__3674\,
            in1 => \N__2246\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U_MD7AndNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MD7LegalizeSB_DFF_LC_5_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U_MD7LegalizeSB_DFFNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5741\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_ROMEN1_NLegalizeSB_DFF_LC_5_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U_ROMEN1_NLegalizeSB_DFFNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5741\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \UMMU_CASEN.i1_2_lut_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3941\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2720\,
            lcout => \D2_6_N_148\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_ROMEN.i2202_4_lut_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__2435\,
            in1 => \N__2299\,
            in2 => \N__2519\,
            in3 => \N__2321\,
            lcout => \ROMEN2_N_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CASEN_N_padLegalizeSB_DFF_LC_8_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CASEN_N_padLegalizeSB_DFFNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5758\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CXXXOUT_padLegalizeSB_DFF_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CXXXOUT_padLegalizeSB_DFFNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5758\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \EN80_N_padLegalizeSB_DFF_LC_8_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \EN80_N_padLegalizeSB_DFFNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5758\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ROMEN2_N_padLegalizeSB_DFF_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ROMEN2_N_padLegalizeSB_DFFNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5758\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_ADDR_DECODER.CXXX_FXXX_I_0_2_lut_3_lut_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__3230\,
            in1 => \N__3160\,
            in2 => \_gnd_net_\,
            in3 => \N__3654\,
            lcout => \DXXX_N_N_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_ADDR_DECODER.CXXX_FXXX_I_0_79_2_lut_3_lut_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__3161\,
            in1 => \_gnd_net_\,
            in2 => \N__3659\,
            in3 => \N__3231\,
            lcout => \FXXX_N_N_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_ADDR_DECODER.i1193_2_lut_3_lut_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__2949\,
            in1 => \N__2317\,
            in2 => \_gnd_net_\,
            in3 => \N__3375\,
            lcout => \D_FXXX\,
            ltout => \D_FXXX_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \UMMU_CASEN.i1_4_lut_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011100000"
        )
    port map (
            in0 => \N__2298\,
            in1 => \N__2597\,
            in2 => \N__2306\,
            in3 => \N__3949\,
            lcout => n966,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_ROMEN.i1_4_lut_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__2962\,
            in1 => \N__2891\,
            in2 => \N__2303\,
            in3 => \N__3378\,
            lcout => \U_MMU_ROMEN.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_ADDR_DECODER.CXXX_I_0_80_2_lut_3_lut_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__3376\,
            in1 => \N__2960\,
            in2 => \_gnd_net_\,
            in3 => \N__5442\,
            lcout => \C8_FXX\,
            ltout => \C8_FXX_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \UMMU_INTERNALS.C8_FXX_I_0_2_lut_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2282\,
            in3 => \N__2671\,
            lcout => \INTC8ACC\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_ROMEN.i1_2_lut_3_lut_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__2672\,
            in1 => \N__3022\,
            in2 => \_gnd_net_\,
            in3 => \N__2708\,
            lcout => \U_MMU_ROMEN.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_ADDR_DECODER.DXXX_N_N_13_I_0_2_lut_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__2961\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3377\,
            lcout => \CXXX\,
            ltout => \CXXX_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_CXXXOUT.i1_4_lut_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__2890\,
            in1 => \N__2492\,
            in2 => \N__2486\,
            in3 => \N__2707\,
            lcout => \CXXXOUT_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_SOFT_SWITCHES_C05X.i2_4_lut_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__2436\,
            in1 => \N__2483\,
            in2 => \N__5612\,
            in3 => \N__2477\,
            lcout => n907,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_ROMEN.i2207_4_lut_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011111111111"
        )
    port map (
            in0 => \N__2511\,
            in1 => \N__2471\,
            in2 => \N__2465\,
            in3 => \N__2438\,
            lcout => \ROMEN1_N_INT\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_ADDR_DECODER.i2172_3_lut_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__2437\,
            in1 => \N__3707\,
            in2 => \_gnd_net_\,
            in3 => \N__2389\,
            lcout => \U_ADDR_DECODER.n2654\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_EN80.i1_3_lut_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__2518\,
            in1 => \N__2356\,
            in2 => \_gnd_net_\,
            in3 => \N__2536\,
            lcout => \EN80_N_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \UMMU_CASEN.i1_2_lut_adj_48_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2357\,
            in2 => \_gnd_net_\,
            in3 => \N__2537\,
            lcout => \CASEN_N_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_SELMB.i2130_3_lut_LC_10_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__5449\,
            in1 => \N__3391\,
            in2 => \_gnd_net_\,
            in3 => \N__4437\,
            lcout => \U_MMU_SELMB.n2610\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_SELMB.i2092_2_lut_LC_10_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3146\,
            in2 => \_gnd_net_\,
            in3 => \N__3211\,
            lcout => \U_MMU_SELMB.n2572\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_SOFT_SWITCHES_C05X.i616_4_lut_LC_10_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__2633\,
            in1 => \N__5537\,
            in2 => \N__5183\,
            in3 => \N__2327\,
            lcout => \HIRES\,
            ltout => \HIRES_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_SELMB.i2_4_lut_LC_10_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000010001"
        )
    port map (
            in0 => \N__2612\,
            in1 => \N__2606\,
            in2 => \N__2600\,
            in3 => \N__3635\,
            lcout => \U_MMU_SELMB.n2516\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_SOFT_SWITCHES_C08X.OUT_FST_ACC_27_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5176\,
            in2 => \_gnd_net_\,
            in3 => \N__3978\,
            lcout => \U_MMU_SOFT_SWITCHES_C08X.OUT_FST_ACC\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU_MMU_SOFT_SWITCHES_C08X.OUT_FST_ACC_27C_net\,
            ce => 'H',
            sr => \N__5593\
        );

    \U_MMU_SOFT_SWITCHES_C08X.WRPROT_28_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011111111111"
        )
    port map (
            in0 => \N__2584\,
            in1 => \N__3980\,
            in2 => \N__2573\,
            in3 => \N__5179\,
            lcout => \WRPROT\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU_MMU_SOFT_SWITCHES_C08X.OUT_FST_ACC_27C_net\,
            ce => 'H',
            sr => \N__5593\
        );

    \U_MMU_SOFT_SWITCHES_C08X.OUT_WREN_32_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101010000000"
        )
    port map (
            in0 => \N__5178\,
            in1 => \N__3979\,
            in2 => \N__2588\,
            in3 => \N__2572\,
            lcout => \U_MMU_SOFT_SWITCHES_C08X.OUT_WREN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU_MMU_SOFT_SWITCHES_C08X.OUT_FST_ACC_27C_net\,
            ce => 'H',
            sr => \N__5593\
        );

    \U_MMU_SOFT_SWITCHES_C08X.RDRAM_26_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__5177\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4935\,
            lcout => \RDRAM\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU_MMU_SOFT_SWITCHES_C08X.OUT_FST_ACC_27C_net\,
            ce => 'H',
            sr => \N__5593\
        );

    \U_SOFT_SWITCHES_C05X.i619_4_lut_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__2642\,
            in1 => \N__2548\,
            in2 => \N__5186\,
            in3 => \N__5595\,
            lcout => \PG2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_ADDR_DECODER.MC0XX_N_I_3_2_lut_3_lut_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__3409\,
            in1 => \N__2948\,
            in2 => \_gnd_net_\,
            in3 => \N__5463\,
            lcout => \U_ADDR_DECODER.MC0XX_N_N_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_SELMB.SELMB_N_I_0_4_lut_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__2561\,
            in1 => \N__3058\,
            in2 => \N__2552\,
            in3 => \N__2768\,
            lcout => \SELMB_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_HOLD_TIME.D_PHI_0_9_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2657\,
            in3 => \_gnd_net_\,
            lcout => \D_PHI_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3296\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \UMMU_INTERNALS.i1172_2_lut_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4239\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2701\,
            lcout => OPEN,
            ltout => \UMMU_INTERNALS.n1605_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \UMMU_INTERNALS.i1_4_lut_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__3005\,
            in1 => \N__5599\,
            in2 => \N__2675\,
            in3 => \N__2670\,
            lcout => \INTC8EN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_HOLD_TIME.SHIFT_REGISTER_i1_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2648\,
            lcout => \U_MMU_HOLD_TIME.SHIFT_REGISTER_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3294\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_HOLD_TIME.SHIFT_REGISTER_i0_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4225\,
            lcout => \U_MMU_HOLD_TIME.SHIFT_REGISTER_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3294\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.i2116_2_lut_3_lut_4_lut_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__4933\,
            in1 => \N__3461\,
            in2 => \N__5390\,
            in3 => \N__4748\,
            lcout => n2596,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_MD7.i1_2_lut_3_lut_4_lut_adj_51_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__3460\,
            in1 => \N__5378\,
            in2 => \N__4940\,
            in3 => \N__4751\,
            lcout => n911,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_MD7.A_3__I_0_26_i2_3_lut_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__2627\,
            in1 => \N__2812\,
            in2 => \_gnd_net_\,
            in3 => \N__5171\,
            lcout => \U_MMU_MD7.n2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_MD7.i2171_2_lut_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2726\,
            in2 => \_gnd_net_\,
            in3 => \N__5172\,
            lcout => OPEN,
            ltout => \U_MMU_MD7.n2658_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_MD7.n2707_bdd_4_lut_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110010011000"
        )
    port map (
            in0 => \N__4749\,
            in1 => \N__2732\,
            in2 => \N__2621\,
            in3 => \N__2618\,
            lcout => \U_MMU_MD7.n2710\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_MD7.A_3__I_0_26_i15_4_lut_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__2759\,
            in1 => \N__2864\,
            in2 => \N__3065\,
            in3 => \N__5391\,
            lcout => \UNGATED_MD7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_MD7.A_c_1_bdd_4_lut_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111110100000"
        )
    port map (
            in0 => \N__3077\,
            in1 => \N__2822\,
            in2 => \N__4759\,
            in3 => \N__4934\,
            lcout => \U_MMU_MD7.n2707\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_SOFT_SWITCHES_C08X.BANK2_30_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5392\,
            lcout => \BANK2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU_MMU_SOFT_SWITCHES_C08X.BANK2_30C_net\,
            ce => 'H',
            sr => \N__5611\
        );

    \U_MMU_SOFT_SWITCHES_C08X.RDROM_31_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4936\,
            in2 => \_gnd_net_\,
            in3 => \N__5105\,
            lcout => \RDROM\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU_MMU_SOFT_SWITCHES_C08X.RDROM_31C_net\,
            ce => 'H',
            sr => \N__5594\
        );

    \U_MMU_SOFT_SWITCHES_C08X.BANK1_25_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5393\,
            lcout => \BANK1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU_MMU_SOFT_SWITCHES_C08X.RDROM_31C_net\,
            ce => 'H',
            sr => \N__5594\
        );

    \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.i631_4_lut_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__2833\,
            in1 => \N__2972\,
            in2 => \N__5607\,
            in3 => \N__5185\,
            lcout => \INTC300_N\,
            ltout => \INTC300_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_ADDR_DECODER.i2_4_lut_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__4448\,
            in1 => \N__3035\,
            in2 => \N__2711\,
            in3 => \N__3106\,
            lcout => \INTC3ACC_N_N_175\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_RA.MMU_RA_MUX.U_DRAM_HOLD_TIME.D_Q3_16_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2870\,
            lcout => \U_MMU_RA.MMU_RA_MUX.D_Q3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_RA.MMU_RA_MUX.U_DRAM_HOLD_TIME.Q3_SHIFT_REGISTER_i0_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4291\,
            lcout => \U_MMU_RA.MMU_RA_MUX.U_DRAM_HOLD_TIME.Q3_SHIFT_REGISTER_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3297\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_RA.MMU_RA_MUX.U_DRAM_HOLD_TIME.Q3_SHIFT_REGISTER_i1_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2876\,
            lcout => \U_MMU_RA.MMU_RA_MUX.U_DRAM_HOLD_TIME.Q3_SHIFT_REGISTER_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3297\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.i2104_2_lut_3_lut_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__5158\,
            in1 => \N__4744\,
            in2 => \_gnd_net_\,
            in3 => \N__4929\,
            lcout => n2584,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.i1_2_lut_4_lut_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__5663\,
            in1 => \N__5309\,
            in2 => \N__4758\,
            in3 => \N__4939\,
            lcout => \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.n2532\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.i614_4_lut_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__5166\,
            in1 => \N__2855\,
            in2 => \N__5606\,
            in3 => \N__2811\,
            lcout => \FLG1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.i1_2_lut_4_lut_4_lut_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__5650\,
            in1 => \N__5339\,
            in2 => \N__4937\,
            in3 => \N__4750\,
            lcout => \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.n937\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.i629_4_lut_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__5591\,
            in1 => \N__5168\,
            in2 => \N__2849\,
            in3 => \N__2794\,
            lcout => \ALTSTKZP\,
            ltout => \ALTSTKZP_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_MD7.A_3__I_0_26_i5_3_lut_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__5167\,
            in1 => \_gnd_net_\,
            in2 => \N__2840\,
            in3 => \N__2837\,
            lcout => \U_MMU_MD7.n5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_ADDR_DECODER.i838_3_lut_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__3950\,
            in1 => \N__5495\,
            in2 => \_gnd_net_\,
            in3 => \N__2816\,
            lcout => OPEN,
            ltout => \SELMB_N_N_137_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_SELMB.SELMB_N_I_24_4_lut_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__2795\,
            in1 => \N__4046\,
            in2 => \N__2783\,
            in3 => \N__2780\,
            lcout => \U_MMU_SELMB.SELMB_N_N_136\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.i1_2_lut_4_lut_adj_50_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__5377\,
            in1 => \N__5664\,
            in2 => \N__4760\,
            in3 => \N__4923\,
            lcout => \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.n938\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_ADDR_DECODER.MA12_I_45_2_lut_3_lut_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__3412\,
            in1 => \N__2966\,
            in2 => \_gnd_net_\,
            in3 => \N__2927\,
            lcout => \MA12_N_209\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_RA.MMU_RA_MUX.U_DRAM_HOLD_TIME.PRAS_N_SHIFT_REGISTER_i0_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4502\,
            lcout => \U_MMU_RA.MMU_RA_MUX.U_DRAM_HOLD_TIME.PRAS_N_SHIFT_REGISTER_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3292\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ORA_pad_6AndLUT4_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2903\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5833\,
            lcout => \ORA_pad_6AndNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ORA_pad_7AndLUT4_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5834\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2897\,
            lcout => \ORA_pad_7AndNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \KBD_N_padLegalizeSB_DFF_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \KBD_N_padLegalizeSB_DFFNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5751\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ORA_pad_6LegalizeSB_DFF_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ORA_pad_6LegalizeSB_DFFNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5751\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ORA_pad_7LegalizeSB_DFF_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ORA_pad_7LegalizeSB_DFFNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5751\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.i1_2_lut_adj_49_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3088\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3821\,
            lcout => \CENROM1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.i633_4_lut_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100010"
        )
    port map (
            in0 => \N__3089\,
            in1 => \N__3836\,
            in2 => \N__5184\,
            in3 => \N__5590\,
            lcout => \PENIO_N\,
            ltout => \PENIO_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_MD7.A_3__I_0_26_i4_3_lut_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5488\,
            in2 => \N__3080\,
            in3 => \N__5162\,
            lcout => \U_MMU_MD7.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.i2090_2_lut_4_lut_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5666\,
            in1 => \N__5376\,
            in2 => \N__4938\,
            in3 => \N__4672\,
            lcout => OPEN,
            ltout => \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.n2570_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.i636_4_lut_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010001010"
        )
    port map (
            in0 => \N__5169\,
            in1 => \N__5592\,
            in2 => \N__3068\,
            in3 => \N__3051\,
            lcout => \EN80VID\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_ADDR_DECODER.i1_2_lut_adj_54_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5239\,
            in2 => \_gnd_net_\,
            in3 => \N__4110\,
            lcout => n927,
            ltout => \n927_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \UMMU_INTERNALS.i2136_4_lut_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3602\,
            in1 => \N__3026\,
            in2 => \N__3011\,
            in3 => \N__3526\,
            lcout => OPEN,
            ltout => \UMMU_INTERNALS.n2616_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \UMMU_INTERNALS.i2142_4_lut_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3434\,
            in1 => \N__3440\,
            in2 => \N__3008\,
            in3 => \N__5170\,
            lcout => \UMMU_INTERNALS.n2622\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_RA.MMU_RA_MUX.COL_RA6_I_0_3_lut_4_lut_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__4592\,
            in1 => \N__4562\,
            in2 => \N__3800\,
            in3 => \N__3236\,
            lcout => \UNGATED_RA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_ADDR_DECODER.i2_3_lut_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__4237\,
            in1 => \N__3703\,
            in2 => \_gnd_net_\,
            in3 => \N__3991\,
            lcout => \KBD_N_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_RA.MMU_RA_MUX.COL_RA7_I_0_3_lut_4_lut_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__4577\,
            in1 => \N__4550\,
            in2 => \N__4115\,
            in3 => \N__3170\,
            lcout => \UNGATED_RA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_RA.MMU_RA_MUX.U_DRAM_HOLD_TIME.PRAS_N_SHIFT_REGISTER_i2_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3242\,
            lcout => \U_MMU_RA.MMU_RA_MUX.U_DRAM_HOLD_TIME.PRAS_N_SHIFT_REGISTER_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3295\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_RA.MMU_RA_MUX.U_DRAM_HOLD_TIME.PRAS_N_SHIFT_REGISTER_i1_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3248\,
            lcout => \U_MMU_RA.MMU_RA_MUX.U_DRAM_HOLD_TIME.PRAS_N_SHIFT_REGISTER_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_MPON.i2_3_lut_4_lut_LC_14_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3650\,
            in1 => \N__4992\,
            in2 => \N__5363\,
            in3 => \N__3229\,
            lcout => \U_MMU_MPON.n2521\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_ADDR_DECODER.i3_4_lut_LC_14_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3649\,
            in1 => \N__3162\,
            in2 => \N__3235\,
            in3 => \N__3410\,
            lcout => \U_ADDR_DECODER.S_0XXX_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_MPON.i2122_4_lut_LC_14_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3592\,
            in1 => \N__5221\,
            in2 => \N__3783\,
            in3 => \N__3163\,
            lcout => OPEN,
            ltout => \U_MMU_MPON.n2602_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_MPON.i2140_4_lut_LC_14_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3411\,
            in1 => \N__3116\,
            in2 => \N__3110\,
            in3 => \N__4430\,
            lcout => n2620,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2096_2_lut_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4232\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3517\,
            lcout => n2576,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_ADDR_DECODER.i2_3_lut_4_lut_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3107\,
            in1 => \N__5232\,
            in2 => \N__4114\,
            in3 => \N__4453\,
            lcout => \MC0XX_N\,
            ltout => \MC0XX_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_ADDR_DECODER.i1_2_lut_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__3788\,
            in1 => \_gnd_net_\,
            in2 => \N__3473\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \n1226_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__3604\,
            in1 => \N__3470\,
            in2 => \N__3464\,
            in3 => \N__4999\,
            lcout => \LATCHED_MC05X_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_MD7.i1_2_lut_adj_52_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4907\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4742\,
            lcout => n933,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \UMMU_INTERNALS.i2100_4_lut_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4236\,
            in1 => \N__3446\,
            in2 => \N__3795\,
            in3 => \N__4447\,
            lcout => \UMMU_INTERNALS.n2580\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_MPON.i1_2_lut_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5000\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5365\,
            lcout => n2520,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_RA.MMU_RA_MUX.D_RAS_N_I_0_2_lut_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__4554\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4591\,
            lcout => OPEN,
            ltout => \U_MMU_RA.MMU_RA_MUX.COMBINED_RAS_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_RA.MMU_RA_MUX.COL_RA4_I_0_4_lut_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__3527\,
            in1 => \N__3428\,
            in2 => \N__3416\,
            in3 => \N__3413\,
            lcout => \UNGATED_RA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_RA.MMU_RA_MUX.U_DRAM_HOLD_TIME.D_RAS_N_14_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3305\,
            lcout => \U_MMU_RA.MMU_RA_MUX.D_RAS_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3298\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_ADDR_DECODER.i293_3_lut_4_lut_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3272\,
            in1 => \N__5459\,
            in2 => \N__5231\,
            in3 => \N__4449\,
            lcout => n626,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_ADDR_DECODER.MMU_1_J5.i2_3_lut_4_lut_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__4982\,
            in1 => \N__3575\,
            in2 => \N__4245\,
            in3 => \N__3510\,
            lcout => n953,
            ltout => \n953_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_DEV_DECODER.MMU_1_P3.i2_3_lut_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111111"
        )
    port map (
            in0 => \N__3826\,
            in1 => \_gnd_net_\,
            in2 => \N__3884\,
            in3 => \N__3761\,
            lcout => \DEV0_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_SOFT_SWITCHES_C00X.i2_3_lut_4_lut_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3992\,
            in1 => \N__3845\,
            in2 => \N__3827\,
            in3 => \N__3787\,
            lcout => \ENABLE_N\,
            ltout => \ENABLE_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_MD7.i1_2_lut_3_lut_4_lut_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__5364\,
            in1 => \N__4713\,
            in2 => \N__3839\,
            in3 => \N__4906\,
            lcout => n912,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_ADDR_DECODER.MMU_1_J5.i1_2_lut_3_lut_4_lut_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3825\,
            in1 => \N__4991\,
            in2 => \N__3799\,
            in3 => \N__3603\,
            lcout => \U_ADDR_DECODER.n44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_ADDR_DECODER.i5_4_lut_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__3896\,
            in1 => \N__4127\,
            in2 => \N__3696\,
            in3 => \N__3525\,
            lcout => \MD7_ENABLE_N_N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_RA.MMU_RA_MUX.COL_RA5_I_0_3_lut_4_lut_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000010"
        )
    port map (
            in0 => \N__3658\,
            in1 => \N__4604\,
            in2 => \N__4561\,
            in3 => \N__3605\,
            lcout => \UNGATED_RA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_MPON.i7_4_lut_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__4016\,
            in1 => \N__4121\,
            in2 => \N__4094\,
            in3 => \N__3524\,
            lcout => n16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_MPON.M5_7_24_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4024\,
            lcout => \U_MMU_MPON.M5_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_ADDR_DECODER.i3_4_lut_adj_53_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011001000"
        )
    port map (
            in0 => \N__3890\,
            in1 => \N__3998\,
            in2 => \N__4246\,
            in3 => \N__5355\,
            lcout => \U_ADDR_DECODER.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_MPON.i4_2_lut_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__4025\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4004\,
            lcout => \U_MMU_MPON.n13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_MPON.M5_2_23_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__4084\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4042\,
            lcout => \U_MMU_MPON.M5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_MPON.DELTA_01XX_N_25_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4015\,
            lcout => \U_MMU_MPON.DELTA_01XX_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_MD7.i2_3_lut_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__4928\,
            in1 => \N__4743\,
            in2 => \_gnd_net_\,
            in3 => \N__5107\,
            lcout => n2523,
            ltout => \n2523_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_ADDR_DECODER.i1_3_lut_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010101010"
        )
    port map (
            in0 => \N__3984\,
            in1 => \_gnd_net_\,
            in2 => \N__3899\,
            in3 => \N__5354\,
            lcout => \U_ADDR_DECODER.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_MD7.i1_2_lut_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4284\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4557\,
            lcout => n906,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_RA.MMU_RA_MUX.i2_3_lut_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__4292\,
            in1 => \N__4501\,
            in2 => \_gnd_net_\,
            in3 => \N__4238\,
            lcout => \U_MMU_RA.MMU_RA_MUX.RA_ENABLE_N_N_215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_RA.MMU_RA_MUX.RA_ENABLE_N_22_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4240\,
            in2 => \_gnd_net_\,
            in3 => \N__4339\,
            lcout => \RA_ENABLE_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU_MMU_RA.MMU_RA_MUX.RA_ENABLE_N_22C_net\,
            ce => 'H',
            sr => \N__4352\
        );

    \RA_ENABLE_N_I_0_1_lut_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4340\,
            lcout => \RA_ENABLE_N_N_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ORA_pad_3AndLUT4_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4310\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5815\,
            lcout => \ORA_pad_3AndNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ORA_pad_4AndLUT4_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5816\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4304\,
            lcout => \ORA_pad_4AndNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ORA_pad_5AndLUT4_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4298\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5817\,
            lcout => \ORA_pad_5AndNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ORA_pad_3LegalizeSB_DFF_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ORA_pad_3LegalizeSB_DFFNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5742\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ORA_pad_4LegalizeSB_DFF_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ORA_pad_4LegalizeSB_DFFNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5742\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ORA_pad_5LegalizeSB_DFF_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ORA_pad_5LegalizeSB_DFFNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5742\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.i1_2_lut_LC_17_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4830\,
            in2 => \_gnd_net_\,
            in3 => \N__4654\,
            lcout => n949,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_MPON.i6_4_lut_LC_17_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__4266\,
            in1 => \N__5465\,
            in2 => \N__4244\,
            in3 => \N__5067\,
            lcout => OPEN,
            ltout => \n15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_SOFT_SWITCHES_C05X.i2199_4_lut_LC_17_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__5693\,
            in1 => \N__5684\,
            in2 => \N__5678\,
            in3 => \N__5675\,
            lcout => \MPON_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.i2086_2_lut_3_lut_4_lut_LC_17_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__5665\,
            in1 => \N__4706\,
            in2 => \N__5313\,
            in3 => \N__4887\,
            lcout => \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.n2566\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_SOFT_SWITCHES_C00X.SOFT_SWITCHES_LATCH.i626_4_lut_LC_17_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__5618\,
            in1 => \N__5527\,
            in2 => \N__5487\,
            in3 => \N__5106\,
            lcout => \FLG2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_RA.MMU_RA_MUX.COL_RA3_I_0_3_lut_4_lut_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__4556\,
            in1 => \N__4617\,
            in2 => \N__5464\,
            in3 => \N__5356\,
            lcout => \UNGATED_RA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_RA.MMU_RA_MUX.COL_RA0_I_0_3_lut_4_lut_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__4616\,
            in1 => \N__4555\,
            in2 => \N__5240\,
            in3 => \N__5157\,
            lcout => \UNGATED_RA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_RA.MMU_RA_MUX.COL_RA1_I_0_3_lut_4_lut_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__4619\,
            in1 => \N__4528\,
            in2 => \N__4970\,
            in3 => \N__4924\,
            lcout => \UNGATED_RA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U_MMU_RA.MMU_RA_MUX.COL_RA2_I_0_3_lut_4_lut_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__4741\,
            in1 => \N__4618\,
            in2 => \N__4549\,
            in3 => \N__4457\,
            lcout => \UNGATED_RA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ORA_pad_0AndLUT4_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5780\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5830\,
            lcout => \ORA_pad_0AndNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ORA_pad_1AndLUT4_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5831\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5774\,
            lcout => \ORA_pad_1AndNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ORA_pad_2AndLUT4_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5768\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5832\,
            lcout => \ORA_pad_2AndNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ORA_pad_0LegalizeSB_DFF_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ORA_pad_0LegalizeSB_DFFNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5732\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ORA_pad_1LegalizeSB_DFF_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ORA_pad_1LegalizeSB_DFFNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5732\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ORA_pad_2LegalizeSB_DFF_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ORA_pad_2LegalizeSB_DFFNet\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5732\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
